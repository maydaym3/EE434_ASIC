module VKSA_128 (in_A, in_B, in_CI, out_S, out_CO);
  input [127:0] in_A, in_B;
  input in_CI;
  output [127:0] out_S;
  output out_CO;

  assign nG_0_0 = in_A[0] & in_B[0];
  assign nP_0_0 = in_A[0] ^ in_B[0];
  assign nG_1_1 = in_A[1] & in_B[1];
  assign nP_1_1 = in_A[1] ^ in_B[1];
  assign nG_2_2 = in_A[2] & in_B[2];
  assign nP_2_2 = in_A[2] ^ in_B[2];
  assign nG_3_3 = in_A[3] & in_B[3];
  assign nP_3_3 = in_A[3] ^ in_B[3];
  assign nG_4_4 = in_A[4] & in_B[4];
  assign nP_4_4 = in_A[4] ^ in_B[4];
  assign nG_5_5 = in_A[5] & in_B[5];
  assign nP_5_5 = in_A[5] ^ in_B[5];
  assign nG_6_6 = in_A[6] & in_B[6];
  assign nP_6_6 = in_A[6] ^ in_B[6];
  assign nG_7_7 = in_A[7] & in_B[7];
  assign nP_7_7 = in_A[7] ^ in_B[7];
  assign nG_8_8 = in_A[8] & in_B[8];
  assign nP_8_8 = in_A[8] ^ in_B[8];
  assign nG_9_9 = in_A[9] & in_B[9];
  assign nP_9_9 = in_A[9] ^ in_B[9];
  assign nG_10_10 = in_A[10] & in_B[10];
  assign nP_10_10 = in_A[10] ^ in_B[10];
  assign nG_11_11 = in_A[11] & in_B[11];
  assign nP_11_11 = in_A[11] ^ in_B[11];
  assign nG_12_12 = in_A[12] & in_B[12];
  assign nP_12_12 = in_A[12] ^ in_B[12];
  assign nG_13_13 = in_A[13] & in_B[13];
  assign nP_13_13 = in_A[13] ^ in_B[13];
  assign nG_14_14 = in_A[14] & in_B[14];
  assign nP_14_14 = in_A[14] ^ in_B[14];
  assign nG_15_15 = in_A[15] & in_B[15];
  assign nP_15_15 = in_A[15] ^ in_B[15];
  assign nG_16_16 = in_A[16] & in_B[16];
  assign nP_16_16 = in_A[16] ^ in_B[16];
  assign nG_17_17 = in_A[17] & in_B[17];
  assign nP_17_17 = in_A[17] ^ in_B[17];
  assign nG_18_18 = in_A[18] & in_B[18];
  assign nP_18_18 = in_A[18] ^ in_B[18];
  assign nG_19_19 = in_A[19] & in_B[19];
  assign nP_19_19 = in_A[19] ^ in_B[19];
  assign nG_20_20 = in_A[20] & in_B[20];
  assign nP_20_20 = in_A[20] ^ in_B[20];
  assign nG_21_21 = in_A[21] & in_B[21];
  assign nP_21_21 = in_A[21] ^ in_B[21];
  assign nG_22_22 = in_A[22] & in_B[22];
  assign nP_22_22 = in_A[22] ^ in_B[22];
  assign nG_23_23 = in_A[23] & in_B[23];
  assign nP_23_23 = in_A[23] ^ in_B[23];
  assign nG_24_24 = in_A[24] & in_B[24];
  assign nP_24_24 = in_A[24] ^ in_B[24];
  assign nG_25_25 = in_A[25] & in_B[25];
  assign nP_25_25 = in_A[25] ^ in_B[25];
  assign nG_26_26 = in_A[26] & in_B[26];
  assign nP_26_26 = in_A[26] ^ in_B[26];
  assign nG_27_27 = in_A[27] & in_B[27];
  assign nP_27_27 = in_A[27] ^ in_B[27];
  assign nG_28_28 = in_A[28] & in_B[28];
  assign nP_28_28 = in_A[28] ^ in_B[28];
  assign nG_29_29 = in_A[29] & in_B[29];
  assign nP_29_29 = in_A[29] ^ in_B[29];
  assign nG_30_30 = in_A[30] & in_B[30];
  assign nP_30_30 = in_A[30] ^ in_B[30];
  assign nG_31_31 = in_A[31] & in_B[31];
  assign nP_31_31 = in_A[31] ^ in_B[31];
  assign nG_32_32 = in_A[32] & in_B[32];
  assign nP_32_32 = in_A[32] ^ in_B[32];
  assign nG_33_33 = in_A[33] & in_B[33];
  assign nP_33_33 = in_A[33] ^ in_B[33];
  assign nG_34_34 = in_A[34] & in_B[34];
  assign nP_34_34 = in_A[34] ^ in_B[34];
  assign nG_35_35 = in_A[35] & in_B[35];
  assign nP_35_35 = in_A[35] ^ in_B[35];
  assign nG_36_36 = in_A[36] & in_B[36];
  assign nP_36_36 = in_A[36] ^ in_B[36];
  assign nG_37_37 = in_A[37] & in_B[37];
  assign nP_37_37 = in_A[37] ^ in_B[37];
  assign nG_38_38 = in_A[38] & in_B[38];
  assign nP_38_38 = in_A[38] ^ in_B[38];
  assign nG_39_39 = in_A[39] & in_B[39];
  assign nP_39_39 = in_A[39] ^ in_B[39];
  assign nG_40_40 = in_A[40] & in_B[40];
  assign nP_40_40 = in_A[40] ^ in_B[40];
  assign nG_41_41 = in_A[41] & in_B[41];
  assign nP_41_41 = in_A[41] ^ in_B[41];
  assign nG_42_42 = in_A[42] & in_B[42];
  assign nP_42_42 = in_A[42] ^ in_B[42];
  assign nG_43_43 = in_A[43] & in_B[43];
  assign nP_43_43 = in_A[43] ^ in_B[43];
  assign nG_44_44 = in_A[44] & in_B[44];
  assign nP_44_44 = in_A[44] ^ in_B[44];
  assign nG_45_45 = in_A[45] & in_B[45];
  assign nP_45_45 = in_A[45] ^ in_B[45];
  assign nG_46_46 = in_A[46] & in_B[46];
  assign nP_46_46 = in_A[46] ^ in_B[46];
  assign nG_47_47 = in_A[47] & in_B[47];
  assign nP_47_47 = in_A[47] ^ in_B[47];
  assign nG_48_48 = in_A[48] & in_B[48];
  assign nP_48_48 = in_A[48] ^ in_B[48];
  assign nG_49_49 = in_A[49] & in_B[49];
  assign nP_49_49 = in_A[49] ^ in_B[49];
  assign nG_50_50 = in_A[50] & in_B[50];
  assign nP_50_50 = in_A[50] ^ in_B[50];
  assign nG_51_51 = in_A[51] & in_B[51];
  assign nP_51_51 = in_A[51] ^ in_B[51];
  assign nG_52_52 = in_A[52] & in_B[52];
  assign nP_52_52 = in_A[52] ^ in_B[52];
  assign nG_53_53 = in_A[53] & in_B[53];
  assign nP_53_53 = in_A[53] ^ in_B[53];
  assign nG_54_54 = in_A[54] & in_B[54];
  assign nP_54_54 = in_A[54] ^ in_B[54];
  assign nG_55_55 = in_A[55] & in_B[55];
  assign nP_55_55 = in_A[55] ^ in_B[55];
  assign nG_56_56 = in_A[56] & in_B[56];
  assign nP_56_56 = in_A[56] ^ in_B[56];
  assign nG_57_57 = in_A[57] & in_B[57];
  assign nP_57_57 = in_A[57] ^ in_B[57];
  assign nG_58_58 = in_A[58] & in_B[58];
  assign nP_58_58 = in_A[58] ^ in_B[58];
  assign nG_59_59 = in_A[59] & in_B[59];
  assign nP_59_59 = in_A[59] ^ in_B[59];
  assign nG_60_60 = in_A[60] & in_B[60];
  assign nP_60_60 = in_A[60] ^ in_B[60];
  assign nG_61_61 = in_A[61] & in_B[61];
  assign nP_61_61 = in_A[61] ^ in_B[61];
  assign nG_62_62 = in_A[62] & in_B[62];
  assign nP_62_62 = in_A[62] ^ in_B[62];
  assign nG_63_63 = in_A[63] & in_B[63];
  assign nP_63_63 = in_A[63] ^ in_B[63];
  assign nG_64_64 = in_A[64] & in_B[64];
  assign nP_64_64 = in_A[64] ^ in_B[64];
  assign nG_65_65 = in_A[65] & in_B[65];
  assign nP_65_65 = in_A[65] ^ in_B[65];
  assign nG_66_66 = in_A[66] & in_B[66];
  assign nP_66_66 = in_A[66] ^ in_B[66];
  assign nG_67_67 = in_A[67] & in_B[67];
  assign nP_67_67 = in_A[67] ^ in_B[67];
  assign nG_68_68 = in_A[68] & in_B[68];
  assign nP_68_68 = in_A[68] ^ in_B[68];
  assign nG_69_69 = in_A[69] & in_B[69];
  assign nP_69_69 = in_A[69] ^ in_B[69];
  assign nG_70_70 = in_A[70] & in_B[70];
  assign nP_70_70 = in_A[70] ^ in_B[70];
  assign nG_71_71 = in_A[71] & in_B[71];
  assign nP_71_71 = in_A[71] ^ in_B[71];
  assign nG_72_72 = in_A[72] & in_B[72];
  assign nP_72_72 = in_A[72] ^ in_B[72];
  assign nG_73_73 = in_A[73] & in_B[73];
  assign nP_73_73 = in_A[73] ^ in_B[73];
  assign nG_74_74 = in_A[74] & in_B[74];
  assign nP_74_74 = in_A[74] ^ in_B[74];
  assign nG_75_75 = in_A[75] & in_B[75];
  assign nP_75_75 = in_A[75] ^ in_B[75];
  assign nG_76_76 = in_A[76] & in_B[76];
  assign nP_76_76 = in_A[76] ^ in_B[76];
  assign nG_77_77 = in_A[77] & in_B[77];
  assign nP_77_77 = in_A[77] ^ in_B[77];
  assign nG_78_78 = in_A[78] & in_B[78];
  assign nP_78_78 = in_A[78] ^ in_B[78];
  assign nG_79_79 = in_A[79] & in_B[79];
  assign nP_79_79 = in_A[79] ^ in_B[79];
  assign nG_80_80 = in_A[80] & in_B[80];
  assign nP_80_80 = in_A[80] ^ in_B[80];
  assign nG_81_81 = in_A[81] & in_B[81];
  assign nP_81_81 = in_A[81] ^ in_B[81];
  assign nG_82_82 = in_A[82] & in_B[82];
  assign nP_82_82 = in_A[82] ^ in_B[82];
  assign nG_83_83 = in_A[83] & in_B[83];
  assign nP_83_83 = in_A[83] ^ in_B[83];
  assign nG_84_84 = in_A[84] & in_B[84];
  assign nP_84_84 = in_A[84] ^ in_B[84];
  assign nG_85_85 = in_A[85] & in_B[85];
  assign nP_85_85 = in_A[85] ^ in_B[85];
  assign nG_86_86 = in_A[86] & in_B[86];
  assign nP_86_86 = in_A[86] ^ in_B[86];
  assign nG_87_87 = in_A[87] & in_B[87];
  assign nP_87_87 = in_A[87] ^ in_B[87];
  assign nG_88_88 = in_A[88] & in_B[88];
  assign nP_88_88 = in_A[88] ^ in_B[88];
  assign nG_89_89 = in_A[89] & in_B[89];
  assign nP_89_89 = in_A[89] ^ in_B[89];
  assign nG_90_90 = in_A[90] & in_B[90];
  assign nP_90_90 = in_A[90] ^ in_B[90];
  assign nG_91_91 = in_A[91] & in_B[91];
  assign nP_91_91 = in_A[91] ^ in_B[91];
  assign nG_92_92 = in_A[92] & in_B[92];
  assign nP_92_92 = in_A[92] ^ in_B[92];
  assign nG_93_93 = in_A[93] & in_B[93];
  assign nP_93_93 = in_A[93] ^ in_B[93];
  assign nG_94_94 = in_A[94] & in_B[94];
  assign nP_94_94 = in_A[94] ^ in_B[94];
  assign nG_95_95 = in_A[95] & in_B[95];
  assign nP_95_95 = in_A[95] ^ in_B[95];
  assign nG_96_96 = in_A[96] & in_B[96];
  assign nP_96_96 = in_A[96] ^ in_B[96];
  assign nG_97_97 = in_A[97] & in_B[97];
  assign nP_97_97 = in_A[97] ^ in_B[97];
  assign nG_98_98 = in_A[98] & in_B[98];
  assign nP_98_98 = in_A[98] ^ in_B[98];
  assign nG_99_99 = in_A[99] & in_B[99];
  assign nP_99_99 = in_A[99] ^ in_B[99];
  assign nG_100_100 = in_A[100] & in_B[100];
  assign nP_100_100 = in_A[100] ^ in_B[100];
  assign nG_101_101 = in_A[101] & in_B[101];
  assign nP_101_101 = in_A[101] ^ in_B[101];
  assign nG_102_102 = in_A[102] & in_B[102];
  assign nP_102_102 = in_A[102] ^ in_B[102];
  assign nG_103_103 = in_A[103] & in_B[103];
  assign nP_103_103 = in_A[103] ^ in_B[103];
  assign nG_104_104 = in_A[104] & in_B[104];
  assign nP_104_104 = in_A[104] ^ in_B[104];
  assign nG_105_105 = in_A[105] & in_B[105];
  assign nP_105_105 = in_A[105] ^ in_B[105];
  assign nG_106_106 = in_A[106] & in_B[106];
  assign nP_106_106 = in_A[106] ^ in_B[106];
  assign nG_107_107 = in_A[107] & in_B[107];
  assign nP_107_107 = in_A[107] ^ in_B[107];
  assign nG_108_108 = in_A[108] & in_B[108];
  assign nP_108_108 = in_A[108] ^ in_B[108];
  assign nG_109_109 = in_A[109] & in_B[109];
  assign nP_109_109 = in_A[109] ^ in_B[109];
  assign nG_110_110 = in_A[110] & in_B[110];
  assign nP_110_110 = in_A[110] ^ in_B[110];
  assign nG_111_111 = in_A[111] & in_B[111];
  assign nP_111_111 = in_A[111] ^ in_B[111];
  assign nG_112_112 = in_A[112] & in_B[112];
  assign nP_112_112 = in_A[112] ^ in_B[112];
  assign nG_113_113 = in_A[113] & in_B[113];
  assign nP_113_113 = in_A[113] ^ in_B[113];
  assign nG_114_114 = in_A[114] & in_B[114];
  assign nP_114_114 = in_A[114] ^ in_B[114];
  assign nG_115_115 = in_A[115] & in_B[115];
  assign nP_115_115 = in_A[115] ^ in_B[115];
  assign nG_116_116 = in_A[116] & in_B[116];
  assign nP_116_116 = in_A[116] ^ in_B[116];
  assign nG_117_117 = in_A[117] & in_B[117];
  assign nP_117_117 = in_A[117] ^ in_B[117];
  assign nG_118_118 = in_A[118] & in_B[118];
  assign nP_118_118 = in_A[118] ^ in_B[118];
  assign nG_119_119 = in_A[119] & in_B[119];
  assign nP_119_119 = in_A[119] ^ in_B[119];
  assign nG_120_120 = in_A[120] & in_B[120];
  assign nP_120_120 = in_A[120] ^ in_B[120];
  assign nG_121_121 = in_A[121] & in_B[121];
  assign nP_121_121 = in_A[121] ^ in_B[121];
  assign nG_122_122 = in_A[122] & in_B[122];
  assign nP_122_122 = in_A[122] ^ in_B[122];
  assign nG_123_123 = in_A[123] & in_B[123];
  assign nP_123_123 = in_A[123] ^ in_B[123];
  assign nG_124_124 = in_A[124] & in_B[124];
  assign nP_124_124 = in_A[124] ^ in_B[124];
  assign nG_125_125 = in_A[125] & in_B[125];
  assign nP_125_125 = in_A[125] ^ in_B[125];
  assign nG_126_126 = in_A[126] & in_B[126];
  assign nP_126_126 = in_A[126] ^ in_B[126];
  assign nG_127_127 = in_A[127] & in_B[127];
  assign nP_127_127 = in_A[127] ^ in_B[127];

  assign nG_127_126 = nG_127_127 | (nP_127_127 & nG_126_126);
  assign nP_127_126 = nP_127_127 & nP_126_126;
  assign nG_126_125 = nG_126_126 | (nP_126_126 & nG_125_125);
  assign nP_126_125 = nP_126_126 & nP_125_125;
  assign nG_125_124 = nG_125_125 | (nP_125_125 & nG_124_124);
  assign nP_125_124 = nP_125_125 & nP_124_124;
  assign nG_124_123 = nG_124_124 | (nP_124_124 & nG_123_123);
  assign nP_124_123 = nP_124_124 & nP_123_123;
  assign nG_123_122 = nG_123_123 | (nP_123_123 & nG_122_122);
  assign nP_123_122 = nP_123_123 & nP_122_122;
  assign nG_122_121 = nG_122_122 | (nP_122_122 & nG_121_121);
  assign nP_122_121 = nP_122_122 & nP_121_121;
  assign nG_121_120 = nG_121_121 | (nP_121_121 & nG_120_120);
  assign nP_121_120 = nP_121_121 & nP_120_120;
  assign nG_120_119 = nG_120_120 | (nP_120_120 & nG_119_119);
  assign nP_120_119 = nP_120_120 & nP_119_119;
  assign nG_119_118 = nG_119_119 | (nP_119_119 & nG_118_118);
  assign nP_119_118 = nP_119_119 & nP_118_118;
  assign nG_118_117 = nG_118_118 | (nP_118_118 & nG_117_117);
  assign nP_118_117 = nP_118_118 & nP_117_117;
  assign nG_117_116 = nG_117_117 | (nP_117_117 & nG_116_116);
  assign nP_117_116 = nP_117_117 & nP_116_116;
  assign nG_116_115 = nG_116_116 | (nP_116_116 & nG_115_115);
  assign nP_116_115 = nP_116_116 & nP_115_115;
  assign nG_115_114 = nG_115_115 | (nP_115_115 & nG_114_114);
  assign nP_115_114 = nP_115_115 & nP_114_114;
  assign nG_114_113 = nG_114_114 | (nP_114_114 & nG_113_113);
  assign nP_114_113 = nP_114_114 & nP_113_113;
  assign nG_113_112 = nG_113_113 | (nP_113_113 & nG_112_112);
  assign nP_113_112 = nP_113_113 & nP_112_112;
  assign nG_112_111 = nG_112_112 | (nP_112_112 & nG_111_111);
  assign nP_112_111 = nP_112_112 & nP_111_111;
  assign nG_111_110 = nG_111_111 | (nP_111_111 & nG_110_110);
  assign nP_111_110 = nP_111_111 & nP_110_110;
  assign nG_110_109 = nG_110_110 | (nP_110_110 & nG_109_109);
  assign nP_110_109 = nP_110_110 & nP_109_109;
  assign nG_109_108 = nG_109_109 | (nP_109_109 & nG_108_108);
  assign nP_109_108 = nP_109_109 & nP_108_108;
  assign nG_108_107 = nG_108_108 | (nP_108_108 & nG_107_107);
  assign nP_108_107 = nP_108_108 & nP_107_107;
  assign nG_107_106 = nG_107_107 | (nP_107_107 & nG_106_106);
  assign nP_107_106 = nP_107_107 & nP_106_106;
  assign nG_106_105 = nG_106_106 | (nP_106_106 & nG_105_105);
  assign nP_106_105 = nP_106_106 & nP_105_105;
  assign nG_105_104 = nG_105_105 | (nP_105_105 & nG_104_104);
  assign nP_105_104 = nP_105_105 & nP_104_104;
  assign nG_104_103 = nG_104_104 | (nP_104_104 & nG_103_103);
  assign nP_104_103 = nP_104_104 & nP_103_103;
  assign nG_103_102 = nG_103_103 | (nP_103_103 & nG_102_102);
  assign nP_103_102 = nP_103_103 & nP_102_102;
  assign nG_102_101 = nG_102_102 | (nP_102_102 & nG_101_101);
  assign nP_102_101 = nP_102_102 & nP_101_101;
  assign nG_101_100 = nG_101_101 | (nP_101_101 & nG_100_100);
  assign nP_101_100 = nP_101_101 & nP_100_100;
  assign nG_100_99 = nG_100_100 | (nP_100_100 & nG_99_99);
  assign nP_100_99 = nP_100_100 & nP_99_99;
  assign nG_99_98 = nG_99_99 | (nP_99_99 & nG_98_98);
  assign nP_99_98 = nP_99_99 & nP_98_98;
  assign nG_98_97 = nG_98_98 | (nP_98_98 & nG_97_97);
  assign nP_98_97 = nP_98_98 & nP_97_97;
  assign nG_97_96 = nG_97_97 | (nP_97_97 & nG_96_96);
  assign nP_97_96 = nP_97_97 & nP_96_96;
  assign nG_96_95 = nG_96_96 | (nP_96_96 & nG_95_95);
  assign nP_96_95 = nP_96_96 & nP_95_95;
  assign nG_95_94 = nG_95_95 | (nP_95_95 & nG_94_94);
  assign nP_95_94 = nP_95_95 & nP_94_94;
  assign nG_94_93 = nG_94_94 | (nP_94_94 & nG_93_93);
  assign nP_94_93 = nP_94_94 & nP_93_93;
  assign nG_93_92 = nG_93_93 | (nP_93_93 & nG_92_92);
  assign nP_93_92 = nP_93_93 & nP_92_92;
  assign nG_92_91 = nG_92_92 | (nP_92_92 & nG_91_91);
  assign nP_92_91 = nP_92_92 & nP_91_91;
  assign nG_91_90 = nG_91_91 | (nP_91_91 & nG_90_90);
  assign nP_91_90 = nP_91_91 & nP_90_90;
  assign nG_90_89 = nG_90_90 | (nP_90_90 & nG_89_89);
  assign nP_90_89 = nP_90_90 & nP_89_89;
  assign nG_89_88 = nG_89_89 | (nP_89_89 & nG_88_88);
  assign nP_89_88 = nP_89_89 & nP_88_88;
  assign nG_88_87 = nG_88_88 | (nP_88_88 & nG_87_87);
  assign nP_88_87 = nP_88_88 & nP_87_87;
  assign nG_87_86 = nG_87_87 | (nP_87_87 & nG_86_86);
  assign nP_87_86 = nP_87_87 & nP_86_86;
  assign nG_86_85 = nG_86_86 | (nP_86_86 & nG_85_85);
  assign nP_86_85 = nP_86_86 & nP_85_85;
  assign nG_85_84 = nG_85_85 | (nP_85_85 & nG_84_84);
  assign nP_85_84 = nP_85_85 & nP_84_84;
  assign nG_84_83 = nG_84_84 | (nP_84_84 & nG_83_83);
  assign nP_84_83 = nP_84_84 & nP_83_83;
  assign nG_83_82 = nG_83_83 | (nP_83_83 & nG_82_82);
  assign nP_83_82 = nP_83_83 & nP_82_82;
  assign nG_82_81 = nG_82_82 | (nP_82_82 & nG_81_81);
  assign nP_82_81 = nP_82_82 & nP_81_81;
  assign nG_81_80 = nG_81_81 | (nP_81_81 & nG_80_80);
  assign nP_81_80 = nP_81_81 & nP_80_80;
  assign nG_80_79 = nG_80_80 | (nP_80_80 & nG_79_79);
  assign nP_80_79 = nP_80_80 & nP_79_79;
  assign nG_79_78 = nG_79_79 | (nP_79_79 & nG_78_78);
  assign nP_79_78 = nP_79_79 & nP_78_78;
  assign nG_78_77 = nG_78_78 | (nP_78_78 & nG_77_77);
  assign nP_78_77 = nP_78_78 & nP_77_77;
  assign nG_77_76 = nG_77_77 | (nP_77_77 & nG_76_76);
  assign nP_77_76 = nP_77_77 & nP_76_76;
  assign nG_76_75 = nG_76_76 | (nP_76_76 & nG_75_75);
  assign nP_76_75 = nP_76_76 & nP_75_75;
  assign nG_75_74 = nG_75_75 | (nP_75_75 & nG_74_74);
  assign nP_75_74 = nP_75_75 & nP_74_74;
  assign nG_74_73 = nG_74_74 | (nP_74_74 & nG_73_73);
  assign nP_74_73 = nP_74_74 & nP_73_73;
  assign nG_73_72 = nG_73_73 | (nP_73_73 & nG_72_72);
  assign nP_73_72 = nP_73_73 & nP_72_72;
  assign nG_72_71 = nG_72_72 | (nP_72_72 & nG_71_71);
  assign nP_72_71 = nP_72_72 & nP_71_71;
  assign nG_71_70 = nG_71_71 | (nP_71_71 & nG_70_70);
  assign nP_71_70 = nP_71_71 & nP_70_70;
  assign nG_70_69 = nG_70_70 | (nP_70_70 & nG_69_69);
  assign nP_70_69 = nP_70_70 & nP_69_69;
  assign nG_69_68 = nG_69_69 | (nP_69_69 & nG_68_68);
  assign nP_69_68 = nP_69_69 & nP_68_68;
  assign nG_68_67 = nG_68_68 | (nP_68_68 & nG_67_67);
  assign nP_68_67 = nP_68_68 & nP_67_67;
  assign nG_67_66 = nG_67_67 | (nP_67_67 & nG_66_66);
  assign nP_67_66 = nP_67_67 & nP_66_66;
  assign nG_66_65 = nG_66_66 | (nP_66_66 & nG_65_65);
  assign nP_66_65 = nP_66_66 & nP_65_65;
  assign nG_65_64 = nG_65_65 | (nP_65_65 & nG_64_64);
  assign nP_65_64 = nP_65_65 & nP_64_64;
  assign nG_64_63 = nG_64_64 | (nP_64_64 & nG_63_63);
  assign nP_64_63 = nP_64_64 & nP_63_63;
  assign nG_63_62 = nG_63_63 | (nP_63_63 & nG_62_62);
  assign nP_63_62 = nP_63_63 & nP_62_62;
  assign nG_62_61 = nG_62_62 | (nP_62_62 & nG_61_61);
  assign nP_62_61 = nP_62_62 & nP_61_61;
  assign nG_61_60 = nG_61_61 | (nP_61_61 & nG_60_60);
  assign nP_61_60 = nP_61_61 & nP_60_60;
  assign nG_60_59 = nG_60_60 | (nP_60_60 & nG_59_59);
  assign nP_60_59 = nP_60_60 & nP_59_59;
  assign nG_59_58 = nG_59_59 | (nP_59_59 & nG_58_58);
  assign nP_59_58 = nP_59_59 & nP_58_58;
  assign nG_58_57 = nG_58_58 | (nP_58_58 & nG_57_57);
  assign nP_58_57 = nP_58_58 & nP_57_57;
  assign nG_57_56 = nG_57_57 | (nP_57_57 & nG_56_56);
  assign nP_57_56 = nP_57_57 & nP_56_56;
  assign nG_56_55 = nG_56_56 | (nP_56_56 & nG_55_55);
  assign nP_56_55 = nP_56_56 & nP_55_55;
  assign nG_55_54 = nG_55_55 | (nP_55_55 & nG_54_54);
  assign nP_55_54 = nP_55_55 & nP_54_54;
  assign nG_54_53 = nG_54_54 | (nP_54_54 & nG_53_53);
  assign nP_54_53 = nP_54_54 & nP_53_53;
  assign nG_53_52 = nG_53_53 | (nP_53_53 & nG_52_52);
  assign nP_53_52 = nP_53_53 & nP_52_52;
  assign nG_52_51 = nG_52_52 | (nP_52_52 & nG_51_51);
  assign nP_52_51 = nP_52_52 & nP_51_51;
  assign nG_51_50 = nG_51_51 | (nP_51_51 & nG_50_50);
  assign nP_51_50 = nP_51_51 & nP_50_50;
  assign nG_50_49 = nG_50_50 | (nP_50_50 & nG_49_49);
  assign nP_50_49 = nP_50_50 & nP_49_49;
  assign nG_49_48 = nG_49_49 | (nP_49_49 & nG_48_48);
  assign nP_49_48 = nP_49_49 & nP_48_48;
  assign nG_48_47 = nG_48_48 | (nP_48_48 & nG_47_47);
  assign nP_48_47 = nP_48_48 & nP_47_47;
  assign nG_47_46 = nG_47_47 | (nP_47_47 & nG_46_46);
  assign nP_47_46 = nP_47_47 & nP_46_46;
  assign nG_46_45 = nG_46_46 | (nP_46_46 & nG_45_45);
  assign nP_46_45 = nP_46_46 & nP_45_45;
  assign nG_45_44 = nG_45_45 | (nP_45_45 & nG_44_44);
  assign nP_45_44 = nP_45_45 & nP_44_44;
  assign nG_44_43 = nG_44_44 | (nP_44_44 & nG_43_43);
  assign nP_44_43 = nP_44_44 & nP_43_43;
  assign nG_43_42 = nG_43_43 | (nP_43_43 & nG_42_42);
  assign nP_43_42 = nP_43_43 & nP_42_42;
  assign nG_42_41 = nG_42_42 | (nP_42_42 & nG_41_41);
  assign nP_42_41 = nP_42_42 & nP_41_41;
  assign nG_41_40 = nG_41_41 | (nP_41_41 & nG_40_40);
  assign nP_41_40 = nP_41_41 & nP_40_40;
  assign nG_40_39 = nG_40_40 | (nP_40_40 & nG_39_39);
  assign nP_40_39 = nP_40_40 & nP_39_39;
  assign nG_39_38 = nG_39_39 | (nP_39_39 & nG_38_38);
  assign nP_39_38 = nP_39_39 & nP_38_38;
  assign nG_38_37 = nG_38_38 | (nP_38_38 & nG_37_37);
  assign nP_38_37 = nP_38_38 & nP_37_37;
  assign nG_37_36 = nG_37_37 | (nP_37_37 & nG_36_36);
  assign nP_37_36 = nP_37_37 & nP_36_36;
  assign nG_36_35 = nG_36_36 | (nP_36_36 & nG_35_35);
  assign nP_36_35 = nP_36_36 & nP_35_35;
  assign nG_35_34 = nG_35_35 | (nP_35_35 & nG_34_34);
  assign nP_35_34 = nP_35_35 & nP_34_34;
  assign nG_34_33 = nG_34_34 | (nP_34_34 & nG_33_33);
  assign nP_34_33 = nP_34_34 & nP_33_33;
  assign nG_33_32 = nG_33_33 | (nP_33_33 & nG_32_32);
  assign nP_33_32 = nP_33_33 & nP_32_32;
  assign nG_32_31 = nG_32_32 | (nP_32_32 & nG_31_31);
  assign nP_32_31 = nP_32_32 & nP_31_31;
  assign nG_31_30 = nG_31_31 | (nP_31_31 & nG_30_30);
  assign nP_31_30 = nP_31_31 & nP_30_30;
  assign nG_30_29 = nG_30_30 | (nP_30_30 & nG_29_29);
  assign nP_30_29 = nP_30_30 & nP_29_29;
  assign nG_29_28 = nG_29_29 | (nP_29_29 & nG_28_28);
  assign nP_29_28 = nP_29_29 & nP_28_28;
  assign nG_28_27 = nG_28_28 | (nP_28_28 & nG_27_27);
  assign nP_28_27 = nP_28_28 & nP_27_27;
  assign nG_27_26 = nG_27_27 | (nP_27_27 & nG_26_26);
  assign nP_27_26 = nP_27_27 & nP_26_26;
  assign nG_26_25 = nG_26_26 | (nP_26_26 & nG_25_25);
  assign nP_26_25 = nP_26_26 & nP_25_25;
  assign nG_25_24 = nG_25_25 | (nP_25_25 & nG_24_24);
  assign nP_25_24 = nP_25_25 & nP_24_24;
  assign nG_24_23 = nG_24_24 | (nP_24_24 & nG_23_23);
  assign nP_24_23 = nP_24_24 & nP_23_23;
  assign nG_23_22 = nG_23_23 | (nP_23_23 & nG_22_22);
  assign nP_23_22 = nP_23_23 & nP_22_22;
  assign nG_22_21 = nG_22_22 | (nP_22_22 & nG_21_21);
  assign nP_22_21 = nP_22_22 & nP_21_21;
  assign nG_21_20 = nG_21_21 | (nP_21_21 & nG_20_20);
  assign nP_21_20 = nP_21_21 & nP_20_20;
  assign nG_20_19 = nG_20_20 | (nP_20_20 & nG_19_19);
  assign nP_20_19 = nP_20_20 & nP_19_19;
  assign nG_19_18 = nG_19_19 | (nP_19_19 & nG_18_18);
  assign nP_19_18 = nP_19_19 & nP_18_18;
  assign nG_18_17 = nG_18_18 | (nP_18_18 & nG_17_17);
  assign nP_18_17 = nP_18_18 & nP_17_17;
  assign nG_17_16 = nG_17_17 | (nP_17_17 & nG_16_16);
  assign nP_17_16 = nP_17_17 & nP_16_16;
  assign nG_16_15 = nG_16_16 | (nP_16_16 & nG_15_15);
  assign nP_16_15 = nP_16_16 & nP_15_15;
  assign nG_15_14 = nG_15_15 | (nP_15_15 & nG_14_14);
  assign nP_15_14 = nP_15_15 & nP_14_14;
  assign nG_14_13 = nG_14_14 | (nP_14_14 & nG_13_13);
  assign nP_14_13 = nP_14_14 & nP_13_13;
  assign nG_13_12 = nG_13_13 | (nP_13_13 & nG_12_12);
  assign nP_13_12 = nP_13_13 & nP_12_12;
  assign nG_12_11 = nG_12_12 | (nP_12_12 & nG_11_11);
  assign nP_12_11 = nP_12_12 & nP_11_11;
  assign nG_11_10 = nG_11_11 | (nP_11_11 & nG_10_10);
  assign nP_11_10 = nP_11_11 & nP_10_10;
  assign nG_10_9 = nG_10_10 | (nP_10_10 & nG_9_9);
  assign nP_10_9 = nP_10_10 & nP_9_9;
  assign nG_9_8 = nG_9_9 | (nP_9_9 & nG_8_8);
  assign nP_9_8 = nP_9_9 & nP_8_8;
  assign nG_8_7 = nG_8_8 | (nP_8_8 & nG_7_7);
  assign nP_8_7 = nP_8_8 & nP_7_7;
  assign nG_7_6 = nG_7_7 | (nP_7_7 & nG_6_6);
  assign nP_7_6 = nP_7_7 & nP_6_6;
  assign nG_6_5 = nG_6_6 | (nP_6_6 & nG_5_5);
  assign nP_6_5 = nP_6_6 & nP_5_5;
  assign nG_5_4 = nG_5_5 | (nP_5_5 & nG_4_4);
  assign nP_5_4 = nP_5_5 & nP_4_4;
  assign nG_4_3 = nG_4_4 | (nP_4_4 & nG_3_3);
  assign nP_4_3 = nP_4_4 & nP_3_3;
  assign nG_3_2 = nG_3_3 | (nP_3_3 & nG_2_2);
  assign nP_3_2 = nP_3_3 & nP_2_2;
  assign nG_2_1 = nG_2_2 | (nP_2_2 & nG_1_1);
  assign nP_2_1 = nP_2_2 & nP_1_1;
  assign nG_1_0 = nG_1_1 | (nP_1_1 & nG_0_0);
  assign nP_1_0 = nP_1_1 & nP_0_0;

  assign nG_127_124 = nG_127_126 | (nP_127_126 & nG_125_124);
  assign nP_127_124 = nP_127_126 & nP_125_124;
  assign nG_126_123 = nG_126_125 | (nP_126_125 & nG_124_123);
  assign nP_126_123 = nP_126_125 & nP_124_123;
  assign nG_125_122 = nG_125_124 | (nP_125_124 & nG_123_122);
  assign nP_125_122 = nP_125_124 & nP_123_122;
  assign nG_124_121 = nG_124_123 | (nP_124_123 & nG_122_121);
  assign nP_124_121 = nP_124_123 & nP_122_121;
  assign nG_123_120 = nG_123_122 | (nP_123_122 & nG_121_120);
  assign nP_123_120 = nP_123_122 & nP_121_120;
  assign nG_122_119 = nG_122_121 | (nP_122_121 & nG_120_119);
  assign nP_122_119 = nP_122_121 & nP_120_119;
  assign nG_121_118 = nG_121_120 | (nP_121_120 & nG_119_118);
  assign nP_121_118 = nP_121_120 & nP_119_118;
  assign nG_120_117 = nG_120_119 | (nP_120_119 & nG_118_117);
  assign nP_120_117 = nP_120_119 & nP_118_117;
  assign nG_119_116 = nG_119_118 | (nP_119_118 & nG_117_116);
  assign nP_119_116 = nP_119_118 & nP_117_116;
  assign nG_118_115 = nG_118_117 | (nP_118_117 & nG_116_115);
  assign nP_118_115 = nP_118_117 & nP_116_115;
  assign nG_117_114 = nG_117_116 | (nP_117_116 & nG_115_114);
  assign nP_117_114 = nP_117_116 & nP_115_114;
  assign nG_116_113 = nG_116_115 | (nP_116_115 & nG_114_113);
  assign nP_116_113 = nP_116_115 & nP_114_113;
  assign nG_115_112 = nG_115_114 | (nP_115_114 & nG_113_112);
  assign nP_115_112 = nP_115_114 & nP_113_112;
  assign nG_114_111 = nG_114_113 | (nP_114_113 & nG_112_111);
  assign nP_114_111 = nP_114_113 & nP_112_111;
  assign nG_113_110 = nG_113_112 | (nP_113_112 & nG_111_110);
  assign nP_113_110 = nP_113_112 & nP_111_110;
  assign nG_112_109 = nG_112_111 | (nP_112_111 & nG_110_109);
  assign nP_112_109 = nP_112_111 & nP_110_109;
  assign nG_111_108 = nG_111_110 | (nP_111_110 & nG_109_108);
  assign nP_111_108 = nP_111_110 & nP_109_108;
  assign nG_110_107 = nG_110_109 | (nP_110_109 & nG_108_107);
  assign nP_110_107 = nP_110_109 & nP_108_107;
  assign nG_109_106 = nG_109_108 | (nP_109_108 & nG_107_106);
  assign nP_109_106 = nP_109_108 & nP_107_106;
  assign nG_108_105 = nG_108_107 | (nP_108_107 & nG_106_105);
  assign nP_108_105 = nP_108_107 & nP_106_105;
  assign nG_107_104 = nG_107_106 | (nP_107_106 & nG_105_104);
  assign nP_107_104 = nP_107_106 & nP_105_104;
  assign nG_106_103 = nG_106_105 | (nP_106_105 & nG_104_103);
  assign nP_106_103 = nP_106_105 & nP_104_103;
  assign nG_105_102 = nG_105_104 | (nP_105_104 & nG_103_102);
  assign nP_105_102 = nP_105_104 & nP_103_102;
  assign nG_104_101 = nG_104_103 | (nP_104_103 & nG_102_101);
  assign nP_104_101 = nP_104_103 & nP_102_101;
  assign nG_103_100 = nG_103_102 | (nP_103_102 & nG_101_100);
  assign nP_103_100 = nP_103_102 & nP_101_100;
  assign nG_102_99 = nG_102_101 | (nP_102_101 & nG_100_99);
  assign nP_102_99 = nP_102_101 & nP_100_99;
  assign nG_101_98 = nG_101_100 | (nP_101_100 & nG_99_98);
  assign nP_101_98 = nP_101_100 & nP_99_98;
  assign nG_100_97 = nG_100_99 | (nP_100_99 & nG_98_97);
  assign nP_100_97 = nP_100_99 & nP_98_97;
  assign nG_99_96 = nG_99_98 | (nP_99_98 & nG_97_96);
  assign nP_99_96 = nP_99_98 & nP_97_96;
  assign nG_98_95 = nG_98_97 | (nP_98_97 & nG_96_95);
  assign nP_98_95 = nP_98_97 & nP_96_95;
  assign nG_97_94 = nG_97_96 | (nP_97_96 & nG_95_94);
  assign nP_97_94 = nP_97_96 & nP_95_94;
  assign nG_96_93 = nG_96_95 | (nP_96_95 & nG_94_93);
  assign nP_96_93 = nP_96_95 & nP_94_93;
  assign nG_95_92 = nG_95_94 | (nP_95_94 & nG_93_92);
  assign nP_95_92 = nP_95_94 & nP_93_92;
  assign nG_94_91 = nG_94_93 | (nP_94_93 & nG_92_91);
  assign nP_94_91 = nP_94_93 & nP_92_91;
  assign nG_93_90 = nG_93_92 | (nP_93_92 & nG_91_90);
  assign nP_93_90 = nP_93_92 & nP_91_90;
  assign nG_92_89 = nG_92_91 | (nP_92_91 & nG_90_89);
  assign nP_92_89 = nP_92_91 & nP_90_89;
  assign nG_91_88 = nG_91_90 | (nP_91_90 & nG_89_88);
  assign nP_91_88 = nP_91_90 & nP_89_88;
  assign nG_90_87 = nG_90_89 | (nP_90_89 & nG_88_87);
  assign nP_90_87 = nP_90_89 & nP_88_87;
  assign nG_89_86 = nG_89_88 | (nP_89_88 & nG_87_86);
  assign nP_89_86 = nP_89_88 & nP_87_86;
  assign nG_88_85 = nG_88_87 | (nP_88_87 & nG_86_85);
  assign nP_88_85 = nP_88_87 & nP_86_85;
  assign nG_87_84 = nG_87_86 | (nP_87_86 & nG_85_84);
  assign nP_87_84 = nP_87_86 & nP_85_84;
  assign nG_86_83 = nG_86_85 | (nP_86_85 & nG_84_83);
  assign nP_86_83 = nP_86_85 & nP_84_83;
  assign nG_85_82 = nG_85_84 | (nP_85_84 & nG_83_82);
  assign nP_85_82 = nP_85_84 & nP_83_82;
  assign nG_84_81 = nG_84_83 | (nP_84_83 & nG_82_81);
  assign nP_84_81 = nP_84_83 & nP_82_81;
  assign nG_83_80 = nG_83_82 | (nP_83_82 & nG_81_80);
  assign nP_83_80 = nP_83_82 & nP_81_80;
  assign nG_82_79 = nG_82_81 | (nP_82_81 & nG_80_79);
  assign nP_82_79 = nP_82_81 & nP_80_79;
  assign nG_81_78 = nG_81_80 | (nP_81_80 & nG_79_78);
  assign nP_81_78 = nP_81_80 & nP_79_78;
  assign nG_80_77 = nG_80_79 | (nP_80_79 & nG_78_77);
  assign nP_80_77 = nP_80_79 & nP_78_77;
  assign nG_79_76 = nG_79_78 | (nP_79_78 & nG_77_76);
  assign nP_79_76 = nP_79_78 & nP_77_76;
  assign nG_78_75 = nG_78_77 | (nP_78_77 & nG_76_75);
  assign nP_78_75 = nP_78_77 & nP_76_75;
  assign nG_77_74 = nG_77_76 | (nP_77_76 & nG_75_74);
  assign nP_77_74 = nP_77_76 & nP_75_74;
  assign nG_76_73 = nG_76_75 | (nP_76_75 & nG_74_73);
  assign nP_76_73 = nP_76_75 & nP_74_73;
  assign nG_75_72 = nG_75_74 | (nP_75_74 & nG_73_72);
  assign nP_75_72 = nP_75_74 & nP_73_72;
  assign nG_74_71 = nG_74_73 | (nP_74_73 & nG_72_71);
  assign nP_74_71 = nP_74_73 & nP_72_71;
  assign nG_73_70 = nG_73_72 | (nP_73_72 & nG_71_70);
  assign nP_73_70 = nP_73_72 & nP_71_70;
  assign nG_72_69 = nG_72_71 | (nP_72_71 & nG_70_69);
  assign nP_72_69 = nP_72_71 & nP_70_69;
  assign nG_71_68 = nG_71_70 | (nP_71_70 & nG_69_68);
  assign nP_71_68 = nP_71_70 & nP_69_68;
  assign nG_70_67 = nG_70_69 | (nP_70_69 & nG_68_67);
  assign nP_70_67 = nP_70_69 & nP_68_67;
  assign nG_69_66 = nG_69_68 | (nP_69_68 & nG_67_66);
  assign nP_69_66 = nP_69_68 & nP_67_66;
  assign nG_68_65 = nG_68_67 | (nP_68_67 & nG_66_65);
  assign nP_68_65 = nP_68_67 & nP_66_65;
  assign nG_67_64 = nG_67_66 | (nP_67_66 & nG_65_64);
  assign nP_67_64 = nP_67_66 & nP_65_64;
  assign nG_66_63 = nG_66_65 | (nP_66_65 & nG_64_63);
  assign nP_66_63 = nP_66_65 & nP_64_63;
  assign nG_65_62 = nG_65_64 | (nP_65_64 & nG_63_62);
  assign nP_65_62 = nP_65_64 & nP_63_62;
  assign nG_64_61 = nG_64_63 | (nP_64_63 & nG_62_61);
  assign nP_64_61 = nP_64_63 & nP_62_61;
  assign nG_63_60 = nG_63_62 | (nP_63_62 & nG_61_60);
  assign nP_63_60 = nP_63_62 & nP_61_60;
  assign nG_62_59 = nG_62_61 | (nP_62_61 & nG_60_59);
  assign nP_62_59 = nP_62_61 & nP_60_59;
  assign nG_61_58 = nG_61_60 | (nP_61_60 & nG_59_58);
  assign nP_61_58 = nP_61_60 & nP_59_58;
  assign nG_60_57 = nG_60_59 | (nP_60_59 & nG_58_57);
  assign nP_60_57 = nP_60_59 & nP_58_57;
  assign nG_59_56 = nG_59_58 | (nP_59_58 & nG_57_56);
  assign nP_59_56 = nP_59_58 & nP_57_56;
  assign nG_58_55 = nG_58_57 | (nP_58_57 & nG_56_55);
  assign nP_58_55 = nP_58_57 & nP_56_55;
  assign nG_57_54 = nG_57_56 | (nP_57_56 & nG_55_54);
  assign nP_57_54 = nP_57_56 & nP_55_54;
  assign nG_56_53 = nG_56_55 | (nP_56_55 & nG_54_53);
  assign nP_56_53 = nP_56_55 & nP_54_53;
  assign nG_55_52 = nG_55_54 | (nP_55_54 & nG_53_52);
  assign nP_55_52 = nP_55_54 & nP_53_52;
  assign nG_54_51 = nG_54_53 | (nP_54_53 & nG_52_51);
  assign nP_54_51 = nP_54_53 & nP_52_51;
  assign nG_53_50 = nG_53_52 | (nP_53_52 & nG_51_50);
  assign nP_53_50 = nP_53_52 & nP_51_50;
  assign nG_52_49 = nG_52_51 | (nP_52_51 & nG_50_49);
  assign nP_52_49 = nP_52_51 & nP_50_49;
  assign nG_51_48 = nG_51_50 | (nP_51_50 & nG_49_48);
  assign nP_51_48 = nP_51_50 & nP_49_48;
  assign nG_50_47 = nG_50_49 | (nP_50_49 & nG_48_47);
  assign nP_50_47 = nP_50_49 & nP_48_47;
  assign nG_49_46 = nG_49_48 | (nP_49_48 & nG_47_46);
  assign nP_49_46 = nP_49_48 & nP_47_46;
  assign nG_48_45 = nG_48_47 | (nP_48_47 & nG_46_45);
  assign nP_48_45 = nP_48_47 & nP_46_45;
  assign nG_47_44 = nG_47_46 | (nP_47_46 & nG_45_44);
  assign nP_47_44 = nP_47_46 & nP_45_44;
  assign nG_46_43 = nG_46_45 | (nP_46_45 & nG_44_43);
  assign nP_46_43 = nP_46_45 & nP_44_43;
  assign nG_45_42 = nG_45_44 | (nP_45_44 & nG_43_42);
  assign nP_45_42 = nP_45_44 & nP_43_42;
  assign nG_44_41 = nG_44_43 | (nP_44_43 & nG_42_41);
  assign nP_44_41 = nP_44_43 & nP_42_41;
  assign nG_43_40 = nG_43_42 | (nP_43_42 & nG_41_40);
  assign nP_43_40 = nP_43_42 & nP_41_40;
  assign nG_42_39 = nG_42_41 | (nP_42_41 & nG_40_39);
  assign nP_42_39 = nP_42_41 & nP_40_39;
  assign nG_41_38 = nG_41_40 | (nP_41_40 & nG_39_38);
  assign nP_41_38 = nP_41_40 & nP_39_38;
  assign nG_40_37 = nG_40_39 | (nP_40_39 & nG_38_37);
  assign nP_40_37 = nP_40_39 & nP_38_37;
  assign nG_39_36 = nG_39_38 | (nP_39_38 & nG_37_36);
  assign nP_39_36 = nP_39_38 & nP_37_36;
  assign nG_38_35 = nG_38_37 | (nP_38_37 & nG_36_35);
  assign nP_38_35 = nP_38_37 & nP_36_35;
  assign nG_37_34 = nG_37_36 | (nP_37_36 & nG_35_34);
  assign nP_37_34 = nP_37_36 & nP_35_34;
  assign nG_36_33 = nG_36_35 | (nP_36_35 & nG_34_33);
  assign nP_36_33 = nP_36_35 & nP_34_33;
  assign nG_35_32 = nG_35_34 | (nP_35_34 & nG_33_32);
  assign nP_35_32 = nP_35_34 & nP_33_32;
  assign nG_34_31 = nG_34_33 | (nP_34_33 & nG_32_31);
  assign nP_34_31 = nP_34_33 & nP_32_31;
  assign nG_33_30 = nG_33_32 | (nP_33_32 & nG_31_30);
  assign nP_33_30 = nP_33_32 & nP_31_30;
  assign nG_32_29 = nG_32_31 | (nP_32_31 & nG_30_29);
  assign nP_32_29 = nP_32_31 & nP_30_29;
  assign nG_31_28 = nG_31_30 | (nP_31_30 & nG_29_28);
  assign nP_31_28 = nP_31_30 & nP_29_28;
  assign nG_30_27 = nG_30_29 | (nP_30_29 & nG_28_27);
  assign nP_30_27 = nP_30_29 & nP_28_27;
  assign nG_29_26 = nG_29_28 | (nP_29_28 & nG_27_26);
  assign nP_29_26 = nP_29_28 & nP_27_26;
  assign nG_28_25 = nG_28_27 | (nP_28_27 & nG_26_25);
  assign nP_28_25 = nP_28_27 & nP_26_25;
  assign nG_27_24 = nG_27_26 | (nP_27_26 & nG_25_24);
  assign nP_27_24 = nP_27_26 & nP_25_24;
  assign nG_26_23 = nG_26_25 | (nP_26_25 & nG_24_23);
  assign nP_26_23 = nP_26_25 & nP_24_23;
  assign nG_25_22 = nG_25_24 | (nP_25_24 & nG_23_22);
  assign nP_25_22 = nP_25_24 & nP_23_22;
  assign nG_24_21 = nG_24_23 | (nP_24_23 & nG_22_21);
  assign nP_24_21 = nP_24_23 & nP_22_21;
  assign nG_23_20 = nG_23_22 | (nP_23_22 & nG_21_20);
  assign nP_23_20 = nP_23_22 & nP_21_20;
  assign nG_22_19 = nG_22_21 | (nP_22_21 & nG_20_19);
  assign nP_22_19 = nP_22_21 & nP_20_19;
  assign nG_21_18 = nG_21_20 | (nP_21_20 & nG_19_18);
  assign nP_21_18 = nP_21_20 & nP_19_18;
  assign nG_20_17 = nG_20_19 | (nP_20_19 & nG_18_17);
  assign nP_20_17 = nP_20_19 & nP_18_17;
  assign nG_19_16 = nG_19_18 | (nP_19_18 & nG_17_16);
  assign nP_19_16 = nP_19_18 & nP_17_16;
  assign nG_18_15 = nG_18_17 | (nP_18_17 & nG_16_15);
  assign nP_18_15 = nP_18_17 & nP_16_15;
  assign nG_17_14 = nG_17_16 | (nP_17_16 & nG_15_14);
  assign nP_17_14 = nP_17_16 & nP_15_14;
  assign nG_16_13 = nG_16_15 | (nP_16_15 & nG_14_13);
  assign nP_16_13 = nP_16_15 & nP_14_13;
  assign nG_15_12 = nG_15_14 | (nP_15_14 & nG_13_12);
  assign nP_15_12 = nP_15_14 & nP_13_12;
  assign nG_14_11 = nG_14_13 | (nP_14_13 & nG_12_11);
  assign nP_14_11 = nP_14_13 & nP_12_11;
  assign nG_13_10 = nG_13_12 | (nP_13_12 & nG_11_10);
  assign nP_13_10 = nP_13_12 & nP_11_10;
  assign nG_12_9 = nG_12_11 | (nP_12_11 & nG_10_9);
  assign nP_12_9 = nP_12_11 & nP_10_9;
  assign nG_11_8 = nG_11_10 | (nP_11_10 & nG_9_8);
  assign nP_11_8 = nP_11_10 & nP_9_8;
  assign nG_10_7 = nG_10_9 | (nP_10_9 & nG_8_7);
  assign nP_10_7 = nP_10_9 & nP_8_7;
  assign nG_9_6 = nG_9_8 | (nP_9_8 & nG_7_6);
  assign nP_9_6 = nP_9_8 & nP_7_6;
  assign nG_8_5 = nG_8_7 | (nP_8_7 & nG_6_5);
  assign nP_8_5 = nP_8_7 & nP_6_5;
  assign nG_7_4 = nG_7_6 | (nP_7_6 & nG_5_4);
  assign nP_7_4 = nP_7_6 & nP_5_4;
  assign nG_6_3 = nG_6_5 | (nP_6_5 & nG_4_3);
  assign nP_6_3 = nP_6_5 & nP_4_3;
  assign nG_5_2 = nG_5_4 | (nP_5_4 & nG_3_2);
  assign nP_5_2 = nP_5_4 & nP_3_2;
  assign nG_4_1 = nG_4_3 | (nP_4_3 & nG_2_1);
  assign nP_4_1 = nP_4_3 & nP_2_1;
  assign nG_3_0 = nG_3_2 | (nP_3_2 & nG_1_0);
  assign nP_3_0 = nP_3_2 & nP_1_0;
  assign nG_2_0 = nG_2_1 | (nP_2_1 & nG_0_0);
  assign nP_2_0 = nP_2_1 & nP_0_0;

  assign nG_127_120 = nG_127_124 | (nP_127_124 & nG_123_120);
  assign nP_127_120 = nP_127_124 & nP_123_120;
  assign nG_126_119 = nG_126_123 | (nP_126_123 & nG_122_119);
  assign nP_126_119 = nP_126_123 & nP_122_119;
  assign nG_125_118 = nG_125_122 | (nP_125_122 & nG_121_118);
  assign nP_125_118 = nP_125_122 & nP_121_118;
  assign nG_124_117 = nG_124_121 | (nP_124_121 & nG_120_117);
  assign nP_124_117 = nP_124_121 & nP_120_117;
  assign nG_123_116 = nG_123_120 | (nP_123_120 & nG_119_116);
  assign nP_123_116 = nP_123_120 & nP_119_116;
  assign nG_122_115 = nG_122_119 | (nP_122_119 & nG_118_115);
  assign nP_122_115 = nP_122_119 & nP_118_115;
  assign nG_121_114 = nG_121_118 | (nP_121_118 & nG_117_114);
  assign nP_121_114 = nP_121_118 & nP_117_114;
  assign nG_120_113 = nG_120_117 | (nP_120_117 & nG_116_113);
  assign nP_120_113 = nP_120_117 & nP_116_113;
  assign nG_119_112 = nG_119_116 | (nP_119_116 & nG_115_112);
  assign nP_119_112 = nP_119_116 & nP_115_112;
  assign nG_118_111 = nG_118_115 | (nP_118_115 & nG_114_111);
  assign nP_118_111 = nP_118_115 & nP_114_111;
  assign nG_117_110 = nG_117_114 | (nP_117_114 & nG_113_110);
  assign nP_117_110 = nP_117_114 & nP_113_110;
  assign nG_116_109 = nG_116_113 | (nP_116_113 & nG_112_109);
  assign nP_116_109 = nP_116_113 & nP_112_109;
  assign nG_115_108 = nG_115_112 | (nP_115_112 & nG_111_108);
  assign nP_115_108 = nP_115_112 & nP_111_108;
  assign nG_114_107 = nG_114_111 | (nP_114_111 & nG_110_107);
  assign nP_114_107 = nP_114_111 & nP_110_107;
  assign nG_113_106 = nG_113_110 | (nP_113_110 & nG_109_106);
  assign nP_113_106 = nP_113_110 & nP_109_106;
  assign nG_112_105 = nG_112_109 | (nP_112_109 & nG_108_105);
  assign nP_112_105 = nP_112_109 & nP_108_105;
  assign nG_111_104 = nG_111_108 | (nP_111_108 & nG_107_104);
  assign nP_111_104 = nP_111_108 & nP_107_104;
  assign nG_110_103 = nG_110_107 | (nP_110_107 & nG_106_103);
  assign nP_110_103 = nP_110_107 & nP_106_103;
  assign nG_109_102 = nG_109_106 | (nP_109_106 & nG_105_102);
  assign nP_109_102 = nP_109_106 & nP_105_102;
  assign nG_108_101 = nG_108_105 | (nP_108_105 & nG_104_101);
  assign nP_108_101 = nP_108_105 & nP_104_101;
  assign nG_107_100 = nG_107_104 | (nP_107_104 & nG_103_100);
  assign nP_107_100 = nP_107_104 & nP_103_100;
  assign nG_106_99 = nG_106_103 | (nP_106_103 & nG_102_99);
  assign nP_106_99 = nP_106_103 & nP_102_99;
  assign nG_105_98 = nG_105_102 | (nP_105_102 & nG_101_98);
  assign nP_105_98 = nP_105_102 & nP_101_98;
  assign nG_104_97 = nG_104_101 | (nP_104_101 & nG_100_97);
  assign nP_104_97 = nP_104_101 & nP_100_97;
  assign nG_103_96 = nG_103_100 | (nP_103_100 & nG_99_96);
  assign nP_103_96 = nP_103_100 & nP_99_96;
  assign nG_102_95 = nG_102_99 | (nP_102_99 & nG_98_95);
  assign nP_102_95 = nP_102_99 & nP_98_95;
  assign nG_101_94 = nG_101_98 | (nP_101_98 & nG_97_94);
  assign nP_101_94 = nP_101_98 & nP_97_94;
  assign nG_100_93 = nG_100_97 | (nP_100_97 & nG_96_93);
  assign nP_100_93 = nP_100_97 & nP_96_93;
  assign nG_99_92 = nG_99_96 | (nP_99_96 & nG_95_92);
  assign nP_99_92 = nP_99_96 & nP_95_92;
  assign nG_98_91 = nG_98_95 | (nP_98_95 & nG_94_91);
  assign nP_98_91 = nP_98_95 & nP_94_91;
  assign nG_97_90 = nG_97_94 | (nP_97_94 & nG_93_90);
  assign nP_97_90 = nP_97_94 & nP_93_90;
  assign nG_96_89 = nG_96_93 | (nP_96_93 & nG_92_89);
  assign nP_96_89 = nP_96_93 & nP_92_89;
  assign nG_95_88 = nG_95_92 | (nP_95_92 & nG_91_88);
  assign nP_95_88 = nP_95_92 & nP_91_88;
  assign nG_94_87 = nG_94_91 | (nP_94_91 & nG_90_87);
  assign nP_94_87 = nP_94_91 & nP_90_87;
  assign nG_93_86 = nG_93_90 | (nP_93_90 & nG_89_86);
  assign nP_93_86 = nP_93_90 & nP_89_86;
  assign nG_92_85 = nG_92_89 | (nP_92_89 & nG_88_85);
  assign nP_92_85 = nP_92_89 & nP_88_85;
  assign nG_91_84 = nG_91_88 | (nP_91_88 & nG_87_84);
  assign nP_91_84 = nP_91_88 & nP_87_84;
  assign nG_90_83 = nG_90_87 | (nP_90_87 & nG_86_83);
  assign nP_90_83 = nP_90_87 & nP_86_83;
  assign nG_89_82 = nG_89_86 | (nP_89_86 & nG_85_82);
  assign nP_89_82 = nP_89_86 & nP_85_82;
  assign nG_88_81 = nG_88_85 | (nP_88_85 & nG_84_81);
  assign nP_88_81 = nP_88_85 & nP_84_81;
  assign nG_87_80 = nG_87_84 | (nP_87_84 & nG_83_80);
  assign nP_87_80 = nP_87_84 & nP_83_80;
  assign nG_86_79 = nG_86_83 | (nP_86_83 & nG_82_79);
  assign nP_86_79 = nP_86_83 & nP_82_79;
  assign nG_85_78 = nG_85_82 | (nP_85_82 & nG_81_78);
  assign nP_85_78 = nP_85_82 & nP_81_78;
  assign nG_84_77 = nG_84_81 | (nP_84_81 & nG_80_77);
  assign nP_84_77 = nP_84_81 & nP_80_77;
  assign nG_83_76 = nG_83_80 | (nP_83_80 & nG_79_76);
  assign nP_83_76 = nP_83_80 & nP_79_76;
  assign nG_82_75 = nG_82_79 | (nP_82_79 & nG_78_75);
  assign nP_82_75 = nP_82_79 & nP_78_75;
  assign nG_81_74 = nG_81_78 | (nP_81_78 & nG_77_74);
  assign nP_81_74 = nP_81_78 & nP_77_74;
  assign nG_80_73 = nG_80_77 | (nP_80_77 & nG_76_73);
  assign nP_80_73 = nP_80_77 & nP_76_73;
  assign nG_79_72 = nG_79_76 | (nP_79_76 & nG_75_72);
  assign nP_79_72 = nP_79_76 & nP_75_72;
  assign nG_78_71 = nG_78_75 | (nP_78_75 & nG_74_71);
  assign nP_78_71 = nP_78_75 & nP_74_71;
  assign nG_77_70 = nG_77_74 | (nP_77_74 & nG_73_70);
  assign nP_77_70 = nP_77_74 & nP_73_70;
  assign nG_76_69 = nG_76_73 | (nP_76_73 & nG_72_69);
  assign nP_76_69 = nP_76_73 & nP_72_69;
  assign nG_75_68 = nG_75_72 | (nP_75_72 & nG_71_68);
  assign nP_75_68 = nP_75_72 & nP_71_68;
  assign nG_74_67 = nG_74_71 | (nP_74_71 & nG_70_67);
  assign nP_74_67 = nP_74_71 & nP_70_67;
  assign nG_73_66 = nG_73_70 | (nP_73_70 & nG_69_66);
  assign nP_73_66 = nP_73_70 & nP_69_66;
  assign nG_72_65 = nG_72_69 | (nP_72_69 & nG_68_65);
  assign nP_72_65 = nP_72_69 & nP_68_65;
  assign nG_71_64 = nG_71_68 | (nP_71_68 & nG_67_64);
  assign nP_71_64 = nP_71_68 & nP_67_64;
  assign nG_70_63 = nG_70_67 | (nP_70_67 & nG_66_63);
  assign nP_70_63 = nP_70_67 & nP_66_63;
  assign nG_69_62 = nG_69_66 | (nP_69_66 & nG_65_62);
  assign nP_69_62 = nP_69_66 & nP_65_62;
  assign nG_68_61 = nG_68_65 | (nP_68_65 & nG_64_61);
  assign nP_68_61 = nP_68_65 & nP_64_61;
  assign nG_67_60 = nG_67_64 | (nP_67_64 & nG_63_60);
  assign nP_67_60 = nP_67_64 & nP_63_60;
  assign nG_66_59 = nG_66_63 | (nP_66_63 & nG_62_59);
  assign nP_66_59 = nP_66_63 & nP_62_59;
  assign nG_65_58 = nG_65_62 | (nP_65_62 & nG_61_58);
  assign nP_65_58 = nP_65_62 & nP_61_58;
  assign nG_64_57 = nG_64_61 | (nP_64_61 & nG_60_57);
  assign nP_64_57 = nP_64_61 & nP_60_57;
  assign nG_63_56 = nG_63_60 | (nP_63_60 & nG_59_56);
  assign nP_63_56 = nP_63_60 & nP_59_56;
  assign nG_62_55 = nG_62_59 | (nP_62_59 & nG_58_55);
  assign nP_62_55 = nP_62_59 & nP_58_55;
  assign nG_61_54 = nG_61_58 | (nP_61_58 & nG_57_54);
  assign nP_61_54 = nP_61_58 & nP_57_54;
  assign nG_60_53 = nG_60_57 | (nP_60_57 & nG_56_53);
  assign nP_60_53 = nP_60_57 & nP_56_53;
  assign nG_59_52 = nG_59_56 | (nP_59_56 & nG_55_52);
  assign nP_59_52 = nP_59_56 & nP_55_52;
  assign nG_58_51 = nG_58_55 | (nP_58_55 & nG_54_51);
  assign nP_58_51 = nP_58_55 & nP_54_51;
  assign nG_57_50 = nG_57_54 | (nP_57_54 & nG_53_50);
  assign nP_57_50 = nP_57_54 & nP_53_50;
  assign nG_56_49 = nG_56_53 | (nP_56_53 & nG_52_49);
  assign nP_56_49 = nP_56_53 & nP_52_49;
  assign nG_55_48 = nG_55_52 | (nP_55_52 & nG_51_48);
  assign nP_55_48 = nP_55_52 & nP_51_48;
  assign nG_54_47 = nG_54_51 | (nP_54_51 & nG_50_47);
  assign nP_54_47 = nP_54_51 & nP_50_47;
  assign nG_53_46 = nG_53_50 | (nP_53_50 & nG_49_46);
  assign nP_53_46 = nP_53_50 & nP_49_46;
  assign nG_52_45 = nG_52_49 | (nP_52_49 & nG_48_45);
  assign nP_52_45 = nP_52_49 & nP_48_45;
  assign nG_51_44 = nG_51_48 | (nP_51_48 & nG_47_44);
  assign nP_51_44 = nP_51_48 & nP_47_44;
  assign nG_50_43 = nG_50_47 | (nP_50_47 & nG_46_43);
  assign nP_50_43 = nP_50_47 & nP_46_43;
  assign nG_49_42 = nG_49_46 | (nP_49_46 & nG_45_42);
  assign nP_49_42 = nP_49_46 & nP_45_42;
  assign nG_48_41 = nG_48_45 | (nP_48_45 & nG_44_41);
  assign nP_48_41 = nP_48_45 & nP_44_41;
  assign nG_47_40 = nG_47_44 | (nP_47_44 & nG_43_40);
  assign nP_47_40 = nP_47_44 & nP_43_40;
  assign nG_46_39 = nG_46_43 | (nP_46_43 & nG_42_39);
  assign nP_46_39 = nP_46_43 & nP_42_39;
  assign nG_45_38 = nG_45_42 | (nP_45_42 & nG_41_38);
  assign nP_45_38 = nP_45_42 & nP_41_38;
  assign nG_44_37 = nG_44_41 | (nP_44_41 & nG_40_37);
  assign nP_44_37 = nP_44_41 & nP_40_37;
  assign nG_43_36 = nG_43_40 | (nP_43_40 & nG_39_36);
  assign nP_43_36 = nP_43_40 & nP_39_36;
  assign nG_42_35 = nG_42_39 | (nP_42_39 & nG_38_35);
  assign nP_42_35 = nP_42_39 & nP_38_35;
  assign nG_41_34 = nG_41_38 | (nP_41_38 & nG_37_34);
  assign nP_41_34 = nP_41_38 & nP_37_34;
  assign nG_40_33 = nG_40_37 | (nP_40_37 & nG_36_33);
  assign nP_40_33 = nP_40_37 & nP_36_33;
  assign nG_39_32 = nG_39_36 | (nP_39_36 & nG_35_32);
  assign nP_39_32 = nP_39_36 & nP_35_32;
  assign nG_38_31 = nG_38_35 | (nP_38_35 & nG_34_31);
  assign nP_38_31 = nP_38_35 & nP_34_31;
  assign nG_37_30 = nG_37_34 | (nP_37_34 & nG_33_30);
  assign nP_37_30 = nP_37_34 & nP_33_30;
  assign nG_36_29 = nG_36_33 | (nP_36_33 & nG_32_29);
  assign nP_36_29 = nP_36_33 & nP_32_29;
  assign nG_35_28 = nG_35_32 | (nP_35_32 & nG_31_28);
  assign nP_35_28 = nP_35_32 & nP_31_28;
  assign nG_34_27 = nG_34_31 | (nP_34_31 & nG_30_27);
  assign nP_34_27 = nP_34_31 & nP_30_27;
  assign nG_33_26 = nG_33_30 | (nP_33_30 & nG_29_26);
  assign nP_33_26 = nP_33_30 & nP_29_26;
  assign nG_32_25 = nG_32_29 | (nP_32_29 & nG_28_25);
  assign nP_32_25 = nP_32_29 & nP_28_25;
  assign nG_31_24 = nG_31_28 | (nP_31_28 & nG_27_24);
  assign nP_31_24 = nP_31_28 & nP_27_24;
  assign nG_30_23 = nG_30_27 | (nP_30_27 & nG_26_23);
  assign nP_30_23 = nP_30_27 & nP_26_23;
  assign nG_29_22 = nG_29_26 | (nP_29_26 & nG_25_22);
  assign nP_29_22 = nP_29_26 & nP_25_22;
  assign nG_28_21 = nG_28_25 | (nP_28_25 & nG_24_21);
  assign nP_28_21 = nP_28_25 & nP_24_21;
  assign nG_27_20 = nG_27_24 | (nP_27_24 & nG_23_20);
  assign nP_27_20 = nP_27_24 & nP_23_20;
  assign nG_26_19 = nG_26_23 | (nP_26_23 & nG_22_19);
  assign nP_26_19 = nP_26_23 & nP_22_19;
  assign nG_25_18 = nG_25_22 | (nP_25_22 & nG_21_18);
  assign nP_25_18 = nP_25_22 & nP_21_18;
  assign nG_24_17 = nG_24_21 | (nP_24_21 & nG_20_17);
  assign nP_24_17 = nP_24_21 & nP_20_17;
  assign nG_23_16 = nG_23_20 | (nP_23_20 & nG_19_16);
  assign nP_23_16 = nP_23_20 & nP_19_16;
  assign nG_22_15 = nG_22_19 | (nP_22_19 & nG_18_15);
  assign nP_22_15 = nP_22_19 & nP_18_15;
  assign nG_21_14 = nG_21_18 | (nP_21_18 & nG_17_14);
  assign nP_21_14 = nP_21_18 & nP_17_14;
  assign nG_20_13 = nG_20_17 | (nP_20_17 & nG_16_13);
  assign nP_20_13 = nP_20_17 & nP_16_13;
  assign nG_19_12 = nG_19_16 | (nP_19_16 & nG_15_12);
  assign nP_19_12 = nP_19_16 & nP_15_12;
  assign nG_18_11 = nG_18_15 | (nP_18_15 & nG_14_11);
  assign nP_18_11 = nP_18_15 & nP_14_11;
  assign nG_17_10 = nG_17_14 | (nP_17_14 & nG_13_10);
  assign nP_17_10 = nP_17_14 & nP_13_10;
  assign nG_16_9 = nG_16_13 | (nP_16_13 & nG_12_9);
  assign nP_16_9 = nP_16_13 & nP_12_9;
  assign nG_15_8 = nG_15_12 | (nP_15_12 & nG_11_8);
  assign nP_15_8 = nP_15_12 & nP_11_8;
  assign nG_14_7 = nG_14_11 | (nP_14_11 & nG_10_7);
  assign nP_14_7 = nP_14_11 & nP_10_7;
  assign nG_13_6 = nG_13_10 | (nP_13_10 & nG_9_6);
  assign nP_13_6 = nP_13_10 & nP_9_6;
  assign nG_12_5 = nG_12_9 | (nP_12_9 & nG_8_5);
  assign nP_12_5 = nP_12_9 & nP_8_5;
  assign nG_11_4 = nG_11_8 | (nP_11_8 & nG_7_4);
  assign nP_11_4 = nP_11_8 & nP_7_4;
  assign nG_10_3 = nG_10_7 | (nP_10_7 & nG_6_3);
  assign nP_10_3 = nP_10_7 & nP_6_3;
  assign nG_9_2 = nG_9_6 | (nP_9_6 & nG_5_2);
  assign nP_9_2 = nP_9_6 & nP_5_2;
  assign nG_8_1 = nG_8_5 | (nP_8_5 & nG_4_1);
  assign nP_8_1 = nP_8_5 & nP_4_1;
  assign nG_7_0 = nG_7_4 | (nP_7_4 & nG_3_0);
  assign nP_7_0 = nP_7_4 & nP_3_0;
  assign nG_6_0 = nG_6_3 | (nP_6_3 & nG_2_0);
  assign nP_6_0 = nP_6_3 & nP_2_0;
  assign nG_5_0 = nG_5_2 | (nP_5_2 & nG_1_0);
  assign nP_5_0 = nP_5_2 & nP_1_0;
  assign nG_4_0 = nG_4_1 | (nP_4_1 & nG_0_0);
  assign nP_4_0 = nP_4_1 & nP_0_0;

  assign nG_127_112 = nG_127_120 | (nP_127_120 & nG_119_112);
  assign nP_127_112 = nP_127_120 & nP_119_112;
  assign nG_126_111 = nG_126_119 | (nP_126_119 & nG_118_111);
  assign nP_126_111 = nP_126_119 & nP_118_111;
  assign nG_125_110 = nG_125_118 | (nP_125_118 & nG_117_110);
  assign nP_125_110 = nP_125_118 & nP_117_110;
  assign nG_124_109 = nG_124_117 | (nP_124_117 & nG_116_109);
  assign nP_124_109 = nP_124_117 & nP_116_109;
  assign nG_123_108 = nG_123_116 | (nP_123_116 & nG_115_108);
  assign nP_123_108 = nP_123_116 & nP_115_108;
  assign nG_122_107 = nG_122_115 | (nP_122_115 & nG_114_107);
  assign nP_122_107 = nP_122_115 & nP_114_107;
  assign nG_121_106 = nG_121_114 | (nP_121_114 & nG_113_106);
  assign nP_121_106 = nP_121_114 & nP_113_106;
  assign nG_120_105 = nG_120_113 | (nP_120_113 & nG_112_105);
  assign nP_120_105 = nP_120_113 & nP_112_105;
  assign nG_119_104 = nG_119_112 | (nP_119_112 & nG_111_104);
  assign nP_119_104 = nP_119_112 & nP_111_104;
  assign nG_118_103 = nG_118_111 | (nP_118_111 & nG_110_103);
  assign nP_118_103 = nP_118_111 & nP_110_103;
  assign nG_117_102 = nG_117_110 | (nP_117_110 & nG_109_102);
  assign nP_117_102 = nP_117_110 & nP_109_102;
  assign nG_116_101 = nG_116_109 | (nP_116_109 & nG_108_101);
  assign nP_116_101 = nP_116_109 & nP_108_101;
  assign nG_115_100 = nG_115_108 | (nP_115_108 & nG_107_100);
  assign nP_115_100 = nP_115_108 & nP_107_100;
  assign nG_114_99 = nG_114_107 | (nP_114_107 & nG_106_99);
  assign nP_114_99 = nP_114_107 & nP_106_99;
  assign nG_113_98 = nG_113_106 | (nP_113_106 & nG_105_98);
  assign nP_113_98 = nP_113_106 & nP_105_98;
  assign nG_112_97 = nG_112_105 | (nP_112_105 & nG_104_97);
  assign nP_112_97 = nP_112_105 & nP_104_97;
  assign nG_111_96 = nG_111_104 | (nP_111_104 & nG_103_96);
  assign nP_111_96 = nP_111_104 & nP_103_96;
  assign nG_110_95 = nG_110_103 | (nP_110_103 & nG_102_95);
  assign nP_110_95 = nP_110_103 & nP_102_95;
  assign nG_109_94 = nG_109_102 | (nP_109_102 & nG_101_94);
  assign nP_109_94 = nP_109_102 & nP_101_94;
  assign nG_108_93 = nG_108_101 | (nP_108_101 & nG_100_93);
  assign nP_108_93 = nP_108_101 & nP_100_93;
  assign nG_107_92 = nG_107_100 | (nP_107_100 & nG_99_92);
  assign nP_107_92 = nP_107_100 & nP_99_92;
  assign nG_106_91 = nG_106_99 | (nP_106_99 & nG_98_91);
  assign nP_106_91 = nP_106_99 & nP_98_91;
  assign nG_105_90 = nG_105_98 | (nP_105_98 & nG_97_90);
  assign nP_105_90 = nP_105_98 & nP_97_90;
  assign nG_104_89 = nG_104_97 | (nP_104_97 & nG_96_89);
  assign nP_104_89 = nP_104_97 & nP_96_89;
  assign nG_103_88 = nG_103_96 | (nP_103_96 & nG_95_88);
  assign nP_103_88 = nP_103_96 & nP_95_88;
  assign nG_102_87 = nG_102_95 | (nP_102_95 & nG_94_87);
  assign nP_102_87 = nP_102_95 & nP_94_87;
  assign nG_101_86 = nG_101_94 | (nP_101_94 & nG_93_86);
  assign nP_101_86 = nP_101_94 & nP_93_86;
  assign nG_100_85 = nG_100_93 | (nP_100_93 & nG_92_85);
  assign nP_100_85 = nP_100_93 & nP_92_85;
  assign nG_99_84 = nG_99_92 | (nP_99_92 & nG_91_84);
  assign nP_99_84 = nP_99_92 & nP_91_84;
  assign nG_98_83 = nG_98_91 | (nP_98_91 & nG_90_83);
  assign nP_98_83 = nP_98_91 & nP_90_83;
  assign nG_97_82 = nG_97_90 | (nP_97_90 & nG_89_82);
  assign nP_97_82 = nP_97_90 & nP_89_82;
  assign nG_96_81 = nG_96_89 | (nP_96_89 & nG_88_81);
  assign nP_96_81 = nP_96_89 & nP_88_81;
  assign nG_95_80 = nG_95_88 | (nP_95_88 & nG_87_80);
  assign nP_95_80 = nP_95_88 & nP_87_80;
  assign nG_94_79 = nG_94_87 | (nP_94_87 & nG_86_79);
  assign nP_94_79 = nP_94_87 & nP_86_79;
  assign nG_93_78 = nG_93_86 | (nP_93_86 & nG_85_78);
  assign nP_93_78 = nP_93_86 & nP_85_78;
  assign nG_92_77 = nG_92_85 | (nP_92_85 & nG_84_77);
  assign nP_92_77 = nP_92_85 & nP_84_77;
  assign nG_91_76 = nG_91_84 | (nP_91_84 & nG_83_76);
  assign nP_91_76 = nP_91_84 & nP_83_76;
  assign nG_90_75 = nG_90_83 | (nP_90_83 & nG_82_75);
  assign nP_90_75 = nP_90_83 & nP_82_75;
  assign nG_89_74 = nG_89_82 | (nP_89_82 & nG_81_74);
  assign nP_89_74 = nP_89_82 & nP_81_74;
  assign nG_88_73 = nG_88_81 | (nP_88_81 & nG_80_73);
  assign nP_88_73 = nP_88_81 & nP_80_73;
  assign nG_87_72 = nG_87_80 | (nP_87_80 & nG_79_72);
  assign nP_87_72 = nP_87_80 & nP_79_72;
  assign nG_86_71 = nG_86_79 | (nP_86_79 & nG_78_71);
  assign nP_86_71 = nP_86_79 & nP_78_71;
  assign nG_85_70 = nG_85_78 | (nP_85_78 & nG_77_70);
  assign nP_85_70 = nP_85_78 & nP_77_70;
  assign nG_84_69 = nG_84_77 | (nP_84_77 & nG_76_69);
  assign nP_84_69 = nP_84_77 & nP_76_69;
  assign nG_83_68 = nG_83_76 | (nP_83_76 & nG_75_68);
  assign nP_83_68 = nP_83_76 & nP_75_68;
  assign nG_82_67 = nG_82_75 | (nP_82_75 & nG_74_67);
  assign nP_82_67 = nP_82_75 & nP_74_67;
  assign nG_81_66 = nG_81_74 | (nP_81_74 & nG_73_66);
  assign nP_81_66 = nP_81_74 & nP_73_66;
  assign nG_80_65 = nG_80_73 | (nP_80_73 & nG_72_65);
  assign nP_80_65 = nP_80_73 & nP_72_65;
  assign nG_79_64 = nG_79_72 | (nP_79_72 & nG_71_64);
  assign nP_79_64 = nP_79_72 & nP_71_64;
  assign nG_78_63 = nG_78_71 | (nP_78_71 & nG_70_63);
  assign nP_78_63 = nP_78_71 & nP_70_63;
  assign nG_77_62 = nG_77_70 | (nP_77_70 & nG_69_62);
  assign nP_77_62 = nP_77_70 & nP_69_62;
  assign nG_76_61 = nG_76_69 | (nP_76_69 & nG_68_61);
  assign nP_76_61 = nP_76_69 & nP_68_61;
  assign nG_75_60 = nG_75_68 | (nP_75_68 & nG_67_60);
  assign nP_75_60 = nP_75_68 & nP_67_60;
  assign nG_74_59 = nG_74_67 | (nP_74_67 & nG_66_59);
  assign nP_74_59 = nP_74_67 & nP_66_59;
  assign nG_73_58 = nG_73_66 | (nP_73_66 & nG_65_58);
  assign nP_73_58 = nP_73_66 & nP_65_58;
  assign nG_72_57 = nG_72_65 | (nP_72_65 & nG_64_57);
  assign nP_72_57 = nP_72_65 & nP_64_57;
  assign nG_71_56 = nG_71_64 | (nP_71_64 & nG_63_56);
  assign nP_71_56 = nP_71_64 & nP_63_56;
  assign nG_70_55 = nG_70_63 | (nP_70_63 & nG_62_55);
  assign nP_70_55 = nP_70_63 & nP_62_55;
  assign nG_69_54 = nG_69_62 | (nP_69_62 & nG_61_54);
  assign nP_69_54 = nP_69_62 & nP_61_54;
  assign nG_68_53 = nG_68_61 | (nP_68_61 & nG_60_53);
  assign nP_68_53 = nP_68_61 & nP_60_53;
  assign nG_67_52 = nG_67_60 | (nP_67_60 & nG_59_52);
  assign nP_67_52 = nP_67_60 & nP_59_52;
  assign nG_66_51 = nG_66_59 | (nP_66_59 & nG_58_51);
  assign nP_66_51 = nP_66_59 & nP_58_51;
  assign nG_65_50 = nG_65_58 | (nP_65_58 & nG_57_50);
  assign nP_65_50 = nP_65_58 & nP_57_50;
  assign nG_64_49 = nG_64_57 | (nP_64_57 & nG_56_49);
  assign nP_64_49 = nP_64_57 & nP_56_49;
  assign nG_63_48 = nG_63_56 | (nP_63_56 & nG_55_48);
  assign nP_63_48 = nP_63_56 & nP_55_48;
  assign nG_62_47 = nG_62_55 | (nP_62_55 & nG_54_47);
  assign nP_62_47 = nP_62_55 & nP_54_47;
  assign nG_61_46 = nG_61_54 | (nP_61_54 & nG_53_46);
  assign nP_61_46 = nP_61_54 & nP_53_46;
  assign nG_60_45 = nG_60_53 | (nP_60_53 & nG_52_45);
  assign nP_60_45 = nP_60_53 & nP_52_45;
  assign nG_59_44 = nG_59_52 | (nP_59_52 & nG_51_44);
  assign nP_59_44 = nP_59_52 & nP_51_44;
  assign nG_58_43 = nG_58_51 | (nP_58_51 & nG_50_43);
  assign nP_58_43 = nP_58_51 & nP_50_43;
  assign nG_57_42 = nG_57_50 | (nP_57_50 & nG_49_42);
  assign nP_57_42 = nP_57_50 & nP_49_42;
  assign nG_56_41 = nG_56_49 | (nP_56_49 & nG_48_41);
  assign nP_56_41 = nP_56_49 & nP_48_41;
  assign nG_55_40 = nG_55_48 | (nP_55_48 & nG_47_40);
  assign nP_55_40 = nP_55_48 & nP_47_40;
  assign nG_54_39 = nG_54_47 | (nP_54_47 & nG_46_39);
  assign nP_54_39 = nP_54_47 & nP_46_39;
  assign nG_53_38 = nG_53_46 | (nP_53_46 & nG_45_38);
  assign nP_53_38 = nP_53_46 & nP_45_38;
  assign nG_52_37 = nG_52_45 | (nP_52_45 & nG_44_37);
  assign nP_52_37 = nP_52_45 & nP_44_37;
  assign nG_51_36 = nG_51_44 | (nP_51_44 & nG_43_36);
  assign nP_51_36 = nP_51_44 & nP_43_36;
  assign nG_50_35 = nG_50_43 | (nP_50_43 & nG_42_35);
  assign nP_50_35 = nP_50_43 & nP_42_35;
  assign nG_49_34 = nG_49_42 | (nP_49_42 & nG_41_34);
  assign nP_49_34 = nP_49_42 & nP_41_34;
  assign nG_48_33 = nG_48_41 | (nP_48_41 & nG_40_33);
  assign nP_48_33 = nP_48_41 & nP_40_33;
  assign nG_47_32 = nG_47_40 | (nP_47_40 & nG_39_32);
  assign nP_47_32 = nP_47_40 & nP_39_32;
  assign nG_46_31 = nG_46_39 | (nP_46_39 & nG_38_31);
  assign nP_46_31 = nP_46_39 & nP_38_31;
  assign nG_45_30 = nG_45_38 | (nP_45_38 & nG_37_30);
  assign nP_45_30 = nP_45_38 & nP_37_30;
  assign nG_44_29 = nG_44_37 | (nP_44_37 & nG_36_29);
  assign nP_44_29 = nP_44_37 & nP_36_29;
  assign nG_43_28 = nG_43_36 | (nP_43_36 & nG_35_28);
  assign nP_43_28 = nP_43_36 & nP_35_28;
  assign nG_42_27 = nG_42_35 | (nP_42_35 & nG_34_27);
  assign nP_42_27 = nP_42_35 & nP_34_27;
  assign nG_41_26 = nG_41_34 | (nP_41_34 & nG_33_26);
  assign nP_41_26 = nP_41_34 & nP_33_26;
  assign nG_40_25 = nG_40_33 | (nP_40_33 & nG_32_25);
  assign nP_40_25 = nP_40_33 & nP_32_25;
  assign nG_39_24 = nG_39_32 | (nP_39_32 & nG_31_24);
  assign nP_39_24 = nP_39_32 & nP_31_24;
  assign nG_38_23 = nG_38_31 | (nP_38_31 & nG_30_23);
  assign nP_38_23 = nP_38_31 & nP_30_23;
  assign nG_37_22 = nG_37_30 | (nP_37_30 & nG_29_22);
  assign nP_37_22 = nP_37_30 & nP_29_22;
  assign nG_36_21 = nG_36_29 | (nP_36_29 & nG_28_21);
  assign nP_36_21 = nP_36_29 & nP_28_21;
  assign nG_35_20 = nG_35_28 | (nP_35_28 & nG_27_20);
  assign nP_35_20 = nP_35_28 & nP_27_20;
  assign nG_34_19 = nG_34_27 | (nP_34_27 & nG_26_19);
  assign nP_34_19 = nP_34_27 & nP_26_19;
  assign nG_33_18 = nG_33_26 | (nP_33_26 & nG_25_18);
  assign nP_33_18 = nP_33_26 & nP_25_18;
  assign nG_32_17 = nG_32_25 | (nP_32_25 & nG_24_17);
  assign nP_32_17 = nP_32_25 & nP_24_17;
  assign nG_31_16 = nG_31_24 | (nP_31_24 & nG_23_16);
  assign nP_31_16 = nP_31_24 & nP_23_16;
  assign nG_30_15 = nG_30_23 | (nP_30_23 & nG_22_15);
  assign nP_30_15 = nP_30_23 & nP_22_15;
  assign nG_29_14 = nG_29_22 | (nP_29_22 & nG_21_14);
  assign nP_29_14 = nP_29_22 & nP_21_14;
  assign nG_28_13 = nG_28_21 | (nP_28_21 & nG_20_13);
  assign nP_28_13 = nP_28_21 & nP_20_13;
  assign nG_27_12 = nG_27_20 | (nP_27_20 & nG_19_12);
  assign nP_27_12 = nP_27_20 & nP_19_12;
  assign nG_26_11 = nG_26_19 | (nP_26_19 & nG_18_11);
  assign nP_26_11 = nP_26_19 & nP_18_11;
  assign nG_25_10 = nG_25_18 | (nP_25_18 & nG_17_10);
  assign nP_25_10 = nP_25_18 & nP_17_10;
  assign nG_24_9 = nG_24_17 | (nP_24_17 & nG_16_9);
  assign nP_24_9 = nP_24_17 & nP_16_9;
  assign nG_23_8 = nG_23_16 | (nP_23_16 & nG_15_8);
  assign nP_23_8 = nP_23_16 & nP_15_8;
  assign nG_22_7 = nG_22_15 | (nP_22_15 & nG_14_7);
  assign nP_22_7 = nP_22_15 & nP_14_7;
  assign nG_21_6 = nG_21_14 | (nP_21_14 & nG_13_6);
  assign nP_21_6 = nP_21_14 & nP_13_6;
  assign nG_20_5 = nG_20_13 | (nP_20_13 & nG_12_5);
  assign nP_20_5 = nP_20_13 & nP_12_5;
  assign nG_19_4 = nG_19_12 | (nP_19_12 & nG_11_4);
  assign nP_19_4 = nP_19_12 & nP_11_4;
  assign nG_18_3 = nG_18_11 | (nP_18_11 & nG_10_3);
  assign nP_18_3 = nP_18_11 & nP_10_3;
  assign nG_17_2 = nG_17_10 | (nP_17_10 & nG_9_2);
  assign nP_17_2 = nP_17_10 & nP_9_2;
  assign nG_16_1 = nG_16_9 | (nP_16_9 & nG_8_1);
  assign nP_16_1 = nP_16_9 & nP_8_1;
  assign nG_15_0 = nG_15_8 | (nP_15_8 & nG_7_0);
  assign nP_15_0 = nP_15_8 & nP_7_0;
  assign nG_14_0 = nG_14_7 | (nP_14_7 & nG_6_0);
  assign nP_14_0 = nP_14_7 & nP_6_0;
  assign nG_13_0 = nG_13_6 | (nP_13_6 & nG_5_0);
  assign nP_13_0 = nP_13_6 & nP_5_0;
  assign nG_12_0 = nG_12_5 | (nP_12_5 & nG_4_0);
  assign nP_12_0 = nP_12_5 & nP_4_0;
  assign nG_11_0 = nG_11_4 | (nP_11_4 & nG_3_0);
  assign nP_11_0 = nP_11_4 & nP_3_0;
  assign nG_10_0 = nG_10_3 | (nP_10_3 & nG_2_0);
  assign nP_10_0 = nP_10_3 & nP_2_0;
  assign nG_9_0 = nG_9_2 | (nP_9_2 & nG_1_0);
  assign nP_9_0 = nP_9_2 & nP_1_0;
  assign nG_8_0 = nG_8_1 | (nP_8_1 & nG_0_0);
  assign nP_8_0 = nP_8_1 & nP_0_0;

  assign nG_127_96 = nG_127_112 | (nP_127_112 & nG_111_96);
  assign nP_127_96 = nP_127_112 & nP_111_96;
  assign nG_126_95 = nG_126_111 | (nP_126_111 & nG_110_95);
  assign nP_126_95 = nP_126_111 & nP_110_95;
  assign nG_125_94 = nG_125_110 | (nP_125_110 & nG_109_94);
  assign nP_125_94 = nP_125_110 & nP_109_94;
  assign nG_124_93 = nG_124_109 | (nP_124_109 & nG_108_93);
  assign nP_124_93 = nP_124_109 & nP_108_93;
  assign nG_123_92 = nG_123_108 | (nP_123_108 & nG_107_92);
  assign nP_123_92 = nP_123_108 & nP_107_92;
  assign nG_122_91 = nG_122_107 | (nP_122_107 & nG_106_91);
  assign nP_122_91 = nP_122_107 & nP_106_91;
  assign nG_121_90 = nG_121_106 | (nP_121_106 & nG_105_90);
  assign nP_121_90 = nP_121_106 & nP_105_90;
  assign nG_120_89 = nG_120_105 | (nP_120_105 & nG_104_89);
  assign nP_120_89 = nP_120_105 & nP_104_89;
  assign nG_119_88 = nG_119_104 | (nP_119_104 & nG_103_88);
  assign nP_119_88 = nP_119_104 & nP_103_88;
  assign nG_118_87 = nG_118_103 | (nP_118_103 & nG_102_87);
  assign nP_118_87 = nP_118_103 & nP_102_87;
  assign nG_117_86 = nG_117_102 | (nP_117_102 & nG_101_86);
  assign nP_117_86 = nP_117_102 & nP_101_86;
  assign nG_116_85 = nG_116_101 | (nP_116_101 & nG_100_85);
  assign nP_116_85 = nP_116_101 & nP_100_85;
  assign nG_115_84 = nG_115_100 | (nP_115_100 & nG_99_84);
  assign nP_115_84 = nP_115_100 & nP_99_84;
  assign nG_114_83 = nG_114_99 | (nP_114_99 & nG_98_83);
  assign nP_114_83 = nP_114_99 & nP_98_83;
  assign nG_113_82 = nG_113_98 | (nP_113_98 & nG_97_82);
  assign nP_113_82 = nP_113_98 & nP_97_82;
  assign nG_112_81 = nG_112_97 | (nP_112_97 & nG_96_81);
  assign nP_112_81 = nP_112_97 & nP_96_81;
  assign nG_111_80 = nG_111_96 | (nP_111_96 & nG_95_80);
  assign nP_111_80 = nP_111_96 & nP_95_80;
  assign nG_110_79 = nG_110_95 | (nP_110_95 & nG_94_79);
  assign nP_110_79 = nP_110_95 & nP_94_79;
  assign nG_109_78 = nG_109_94 | (nP_109_94 & nG_93_78);
  assign nP_109_78 = nP_109_94 & nP_93_78;
  assign nG_108_77 = nG_108_93 | (nP_108_93 & nG_92_77);
  assign nP_108_77 = nP_108_93 & nP_92_77;
  assign nG_107_76 = nG_107_92 | (nP_107_92 & nG_91_76);
  assign nP_107_76 = nP_107_92 & nP_91_76;
  assign nG_106_75 = nG_106_91 | (nP_106_91 & nG_90_75);
  assign nP_106_75 = nP_106_91 & nP_90_75;
  assign nG_105_74 = nG_105_90 | (nP_105_90 & nG_89_74);
  assign nP_105_74 = nP_105_90 & nP_89_74;
  assign nG_104_73 = nG_104_89 | (nP_104_89 & nG_88_73);
  assign nP_104_73 = nP_104_89 & nP_88_73;
  assign nG_103_72 = nG_103_88 | (nP_103_88 & nG_87_72);
  assign nP_103_72 = nP_103_88 & nP_87_72;
  assign nG_102_71 = nG_102_87 | (nP_102_87 & nG_86_71);
  assign nP_102_71 = nP_102_87 & nP_86_71;
  assign nG_101_70 = nG_101_86 | (nP_101_86 & nG_85_70);
  assign nP_101_70 = nP_101_86 & nP_85_70;
  assign nG_100_69 = nG_100_85 | (nP_100_85 & nG_84_69);
  assign nP_100_69 = nP_100_85 & nP_84_69;
  assign nG_99_68 = nG_99_84 | (nP_99_84 & nG_83_68);
  assign nP_99_68 = nP_99_84 & nP_83_68;
  assign nG_98_67 = nG_98_83 | (nP_98_83 & nG_82_67);
  assign nP_98_67 = nP_98_83 & nP_82_67;
  assign nG_97_66 = nG_97_82 | (nP_97_82 & nG_81_66);
  assign nP_97_66 = nP_97_82 & nP_81_66;
  assign nG_96_65 = nG_96_81 | (nP_96_81 & nG_80_65);
  assign nP_96_65 = nP_96_81 & nP_80_65;
  assign nG_95_64 = nG_95_80 | (nP_95_80 & nG_79_64);
  assign nP_95_64 = nP_95_80 & nP_79_64;
  assign nG_94_63 = nG_94_79 | (nP_94_79 & nG_78_63);
  assign nP_94_63 = nP_94_79 & nP_78_63;
  assign nG_93_62 = nG_93_78 | (nP_93_78 & nG_77_62);
  assign nP_93_62 = nP_93_78 & nP_77_62;
  assign nG_92_61 = nG_92_77 | (nP_92_77 & nG_76_61);
  assign nP_92_61 = nP_92_77 & nP_76_61;
  assign nG_91_60 = nG_91_76 | (nP_91_76 & nG_75_60);
  assign nP_91_60 = nP_91_76 & nP_75_60;
  assign nG_90_59 = nG_90_75 | (nP_90_75 & nG_74_59);
  assign nP_90_59 = nP_90_75 & nP_74_59;
  assign nG_89_58 = nG_89_74 | (nP_89_74 & nG_73_58);
  assign nP_89_58 = nP_89_74 & nP_73_58;
  assign nG_88_57 = nG_88_73 | (nP_88_73 & nG_72_57);
  assign nP_88_57 = nP_88_73 & nP_72_57;
  assign nG_87_56 = nG_87_72 | (nP_87_72 & nG_71_56);
  assign nP_87_56 = nP_87_72 & nP_71_56;
  assign nG_86_55 = nG_86_71 | (nP_86_71 & nG_70_55);
  assign nP_86_55 = nP_86_71 & nP_70_55;
  assign nG_85_54 = nG_85_70 | (nP_85_70 & nG_69_54);
  assign nP_85_54 = nP_85_70 & nP_69_54;
  assign nG_84_53 = nG_84_69 | (nP_84_69 & nG_68_53);
  assign nP_84_53 = nP_84_69 & nP_68_53;
  assign nG_83_52 = nG_83_68 | (nP_83_68 & nG_67_52);
  assign nP_83_52 = nP_83_68 & nP_67_52;
  assign nG_82_51 = nG_82_67 | (nP_82_67 & nG_66_51);
  assign nP_82_51 = nP_82_67 & nP_66_51;
  assign nG_81_50 = nG_81_66 | (nP_81_66 & nG_65_50);
  assign nP_81_50 = nP_81_66 & nP_65_50;
  assign nG_80_49 = nG_80_65 | (nP_80_65 & nG_64_49);
  assign nP_80_49 = nP_80_65 & nP_64_49;
  assign nG_79_48 = nG_79_64 | (nP_79_64 & nG_63_48);
  assign nP_79_48 = nP_79_64 & nP_63_48;
  assign nG_78_47 = nG_78_63 | (nP_78_63 & nG_62_47);
  assign nP_78_47 = nP_78_63 & nP_62_47;
  assign nG_77_46 = nG_77_62 | (nP_77_62 & nG_61_46);
  assign nP_77_46 = nP_77_62 & nP_61_46;
  assign nG_76_45 = nG_76_61 | (nP_76_61 & nG_60_45);
  assign nP_76_45 = nP_76_61 & nP_60_45;
  assign nG_75_44 = nG_75_60 | (nP_75_60 & nG_59_44);
  assign nP_75_44 = nP_75_60 & nP_59_44;
  assign nG_74_43 = nG_74_59 | (nP_74_59 & nG_58_43);
  assign nP_74_43 = nP_74_59 & nP_58_43;
  assign nG_73_42 = nG_73_58 | (nP_73_58 & nG_57_42);
  assign nP_73_42 = nP_73_58 & nP_57_42;
  assign nG_72_41 = nG_72_57 | (nP_72_57 & nG_56_41);
  assign nP_72_41 = nP_72_57 & nP_56_41;
  assign nG_71_40 = nG_71_56 | (nP_71_56 & nG_55_40);
  assign nP_71_40 = nP_71_56 & nP_55_40;
  assign nG_70_39 = nG_70_55 | (nP_70_55 & nG_54_39);
  assign nP_70_39 = nP_70_55 & nP_54_39;
  assign nG_69_38 = nG_69_54 | (nP_69_54 & nG_53_38);
  assign nP_69_38 = nP_69_54 & nP_53_38;
  assign nG_68_37 = nG_68_53 | (nP_68_53 & nG_52_37);
  assign nP_68_37 = nP_68_53 & nP_52_37;
  assign nG_67_36 = nG_67_52 | (nP_67_52 & nG_51_36);
  assign nP_67_36 = nP_67_52 & nP_51_36;
  assign nG_66_35 = nG_66_51 | (nP_66_51 & nG_50_35);
  assign nP_66_35 = nP_66_51 & nP_50_35;
  assign nG_65_34 = nG_65_50 | (nP_65_50 & nG_49_34);
  assign nP_65_34 = nP_65_50 & nP_49_34;
  assign nG_64_33 = nG_64_49 | (nP_64_49 & nG_48_33);
  assign nP_64_33 = nP_64_49 & nP_48_33;
  assign nG_63_32 = nG_63_48 | (nP_63_48 & nG_47_32);
  assign nP_63_32 = nP_63_48 & nP_47_32;
  assign nG_62_31 = nG_62_47 | (nP_62_47 & nG_46_31);
  assign nP_62_31 = nP_62_47 & nP_46_31;
  assign nG_61_30 = nG_61_46 | (nP_61_46 & nG_45_30);
  assign nP_61_30 = nP_61_46 & nP_45_30;
  assign nG_60_29 = nG_60_45 | (nP_60_45 & nG_44_29);
  assign nP_60_29 = nP_60_45 & nP_44_29;
  assign nG_59_28 = nG_59_44 | (nP_59_44 & nG_43_28);
  assign nP_59_28 = nP_59_44 & nP_43_28;
  assign nG_58_27 = nG_58_43 | (nP_58_43 & nG_42_27);
  assign nP_58_27 = nP_58_43 & nP_42_27;
  assign nG_57_26 = nG_57_42 | (nP_57_42 & nG_41_26);
  assign nP_57_26 = nP_57_42 & nP_41_26;
  assign nG_56_25 = nG_56_41 | (nP_56_41 & nG_40_25);
  assign nP_56_25 = nP_56_41 & nP_40_25;
  assign nG_55_24 = nG_55_40 | (nP_55_40 & nG_39_24);
  assign nP_55_24 = nP_55_40 & nP_39_24;
  assign nG_54_23 = nG_54_39 | (nP_54_39 & nG_38_23);
  assign nP_54_23 = nP_54_39 & nP_38_23;
  assign nG_53_22 = nG_53_38 | (nP_53_38 & nG_37_22);
  assign nP_53_22 = nP_53_38 & nP_37_22;
  assign nG_52_21 = nG_52_37 | (nP_52_37 & nG_36_21);
  assign nP_52_21 = nP_52_37 & nP_36_21;
  assign nG_51_20 = nG_51_36 | (nP_51_36 & nG_35_20);
  assign nP_51_20 = nP_51_36 & nP_35_20;
  assign nG_50_19 = nG_50_35 | (nP_50_35 & nG_34_19);
  assign nP_50_19 = nP_50_35 & nP_34_19;
  assign nG_49_18 = nG_49_34 | (nP_49_34 & nG_33_18);
  assign nP_49_18 = nP_49_34 & nP_33_18;
  assign nG_48_17 = nG_48_33 | (nP_48_33 & nG_32_17);
  assign nP_48_17 = nP_48_33 & nP_32_17;
  assign nG_47_16 = nG_47_32 | (nP_47_32 & nG_31_16);
  assign nP_47_16 = nP_47_32 & nP_31_16;
  assign nG_46_15 = nG_46_31 | (nP_46_31 & nG_30_15);
  assign nP_46_15 = nP_46_31 & nP_30_15;
  assign nG_45_14 = nG_45_30 | (nP_45_30 & nG_29_14);
  assign nP_45_14 = nP_45_30 & nP_29_14;
  assign nG_44_13 = nG_44_29 | (nP_44_29 & nG_28_13);
  assign nP_44_13 = nP_44_29 & nP_28_13;
  assign nG_43_12 = nG_43_28 | (nP_43_28 & nG_27_12);
  assign nP_43_12 = nP_43_28 & nP_27_12;
  assign nG_42_11 = nG_42_27 | (nP_42_27 & nG_26_11);
  assign nP_42_11 = nP_42_27 & nP_26_11;
  assign nG_41_10 = nG_41_26 | (nP_41_26 & nG_25_10);
  assign nP_41_10 = nP_41_26 & nP_25_10;
  assign nG_40_9 = nG_40_25 | (nP_40_25 & nG_24_9);
  assign nP_40_9 = nP_40_25 & nP_24_9;
  assign nG_39_8 = nG_39_24 | (nP_39_24 & nG_23_8);
  assign nP_39_8 = nP_39_24 & nP_23_8;
  assign nG_38_7 = nG_38_23 | (nP_38_23 & nG_22_7);
  assign nP_38_7 = nP_38_23 & nP_22_7;
  assign nG_37_6 = nG_37_22 | (nP_37_22 & nG_21_6);
  assign nP_37_6 = nP_37_22 & nP_21_6;
  assign nG_36_5 = nG_36_21 | (nP_36_21 & nG_20_5);
  assign nP_36_5 = nP_36_21 & nP_20_5;
  assign nG_35_4 = nG_35_20 | (nP_35_20 & nG_19_4);
  assign nP_35_4 = nP_35_20 & nP_19_4;
  assign nG_34_3 = nG_34_19 | (nP_34_19 & nG_18_3);
  assign nP_34_3 = nP_34_19 & nP_18_3;
  assign nG_33_2 = nG_33_18 | (nP_33_18 & nG_17_2);
  assign nP_33_2 = nP_33_18 & nP_17_2;
  assign nG_32_1 = nG_32_17 | (nP_32_17 & nG_16_1);
  assign nP_32_1 = nP_32_17 & nP_16_1;
  assign nG_31_0 = nG_31_16 | (nP_31_16 & nG_15_0);
  assign nP_31_0 = nP_31_16 & nP_15_0;
  assign nG_30_0 = nG_30_15 | (nP_30_15 & nG_14_0);
  assign nP_30_0 = nP_30_15 & nP_14_0;
  assign nG_29_0 = nG_29_14 | (nP_29_14 & nG_13_0);
  assign nP_29_0 = nP_29_14 & nP_13_0;
  assign nG_28_0 = nG_28_13 | (nP_28_13 & nG_12_0);
  assign nP_28_0 = nP_28_13 & nP_12_0;
  assign nG_27_0 = nG_27_12 | (nP_27_12 & nG_11_0);
  assign nP_27_0 = nP_27_12 & nP_11_0;
  assign nG_26_0 = nG_26_11 | (nP_26_11 & nG_10_0);
  assign nP_26_0 = nP_26_11 & nP_10_0;
  assign nG_25_0 = nG_25_10 | (nP_25_10 & nG_9_0);
  assign nP_25_0 = nP_25_10 & nP_9_0;
  assign nG_24_0 = nG_24_9 | (nP_24_9 & nG_8_0);
  assign nP_24_0 = nP_24_9 & nP_8_0;
  assign nG_23_0 = nG_23_8 | (nP_23_8 & nG_7_0);
  assign nP_23_0 = nP_23_8 & nP_7_0;
  assign nG_22_0 = nG_22_7 | (nP_22_7 & nG_6_0);
  assign nP_22_0 = nP_22_7 & nP_6_0;
  assign nG_21_0 = nG_21_6 | (nP_21_6 & nG_5_0);
  assign nP_21_0 = nP_21_6 & nP_5_0;
  assign nG_20_0 = nG_20_5 | (nP_20_5 & nG_4_0);
  assign nP_20_0 = nP_20_5 & nP_4_0;
  assign nG_19_0 = nG_19_4 | (nP_19_4 & nG_3_0);
  assign nP_19_0 = nP_19_4 & nP_3_0;
  assign nG_18_0 = nG_18_3 | (nP_18_3 & nG_2_0);
  assign nP_18_0 = nP_18_3 & nP_2_0;
  assign nG_17_0 = nG_17_2 | (nP_17_2 & nG_1_0);
  assign nP_17_0 = nP_17_2 & nP_1_0;
  assign nG_16_0 = nG_16_1 | (nP_16_1 & nG_0_0);
  assign nP_16_0 = nP_16_1 & nP_0_0;

  assign nG_127_64 = nG_127_96 | (nP_127_96 & nG_95_64);
  assign nP_127_64 = nP_127_96 & nP_95_64;
  assign nG_126_63 = nG_126_95 | (nP_126_95 & nG_94_63);
  assign nP_126_63 = nP_126_95 & nP_94_63;
  assign nG_125_62 = nG_125_94 | (nP_125_94 & nG_93_62);
  assign nP_125_62 = nP_125_94 & nP_93_62;
  assign nG_124_61 = nG_124_93 | (nP_124_93 & nG_92_61);
  assign nP_124_61 = nP_124_93 & nP_92_61;
  assign nG_123_60 = nG_123_92 | (nP_123_92 & nG_91_60);
  assign nP_123_60 = nP_123_92 & nP_91_60;
  assign nG_122_59 = nG_122_91 | (nP_122_91 & nG_90_59);
  assign nP_122_59 = nP_122_91 & nP_90_59;
  assign nG_121_58 = nG_121_90 | (nP_121_90 & nG_89_58);
  assign nP_121_58 = nP_121_90 & nP_89_58;
  assign nG_120_57 = nG_120_89 | (nP_120_89 & nG_88_57);
  assign nP_120_57 = nP_120_89 & nP_88_57;
  assign nG_119_56 = nG_119_88 | (nP_119_88 & nG_87_56);
  assign nP_119_56 = nP_119_88 & nP_87_56;
  assign nG_118_55 = nG_118_87 | (nP_118_87 & nG_86_55);
  assign nP_118_55 = nP_118_87 & nP_86_55;
  assign nG_117_54 = nG_117_86 | (nP_117_86 & nG_85_54);
  assign nP_117_54 = nP_117_86 & nP_85_54;
  assign nG_116_53 = nG_116_85 | (nP_116_85 & nG_84_53);
  assign nP_116_53 = nP_116_85 & nP_84_53;
  assign nG_115_52 = nG_115_84 | (nP_115_84 & nG_83_52);
  assign nP_115_52 = nP_115_84 & nP_83_52;
  assign nG_114_51 = nG_114_83 | (nP_114_83 & nG_82_51);
  assign nP_114_51 = nP_114_83 & nP_82_51;
  assign nG_113_50 = nG_113_82 | (nP_113_82 & nG_81_50);
  assign nP_113_50 = nP_113_82 & nP_81_50;
  assign nG_112_49 = nG_112_81 | (nP_112_81 & nG_80_49);
  assign nP_112_49 = nP_112_81 & nP_80_49;
  assign nG_111_48 = nG_111_80 | (nP_111_80 & nG_79_48);
  assign nP_111_48 = nP_111_80 & nP_79_48;
  assign nG_110_47 = nG_110_79 | (nP_110_79 & nG_78_47);
  assign nP_110_47 = nP_110_79 & nP_78_47;
  assign nG_109_46 = nG_109_78 | (nP_109_78 & nG_77_46);
  assign nP_109_46 = nP_109_78 & nP_77_46;
  assign nG_108_45 = nG_108_77 | (nP_108_77 & nG_76_45);
  assign nP_108_45 = nP_108_77 & nP_76_45;
  assign nG_107_44 = nG_107_76 | (nP_107_76 & nG_75_44);
  assign nP_107_44 = nP_107_76 & nP_75_44;
  assign nG_106_43 = nG_106_75 | (nP_106_75 & nG_74_43);
  assign nP_106_43 = nP_106_75 & nP_74_43;
  assign nG_105_42 = nG_105_74 | (nP_105_74 & nG_73_42);
  assign nP_105_42 = nP_105_74 & nP_73_42;
  assign nG_104_41 = nG_104_73 | (nP_104_73 & nG_72_41);
  assign nP_104_41 = nP_104_73 & nP_72_41;
  assign nG_103_40 = nG_103_72 | (nP_103_72 & nG_71_40);
  assign nP_103_40 = nP_103_72 & nP_71_40;
  assign nG_102_39 = nG_102_71 | (nP_102_71 & nG_70_39);
  assign nP_102_39 = nP_102_71 & nP_70_39;
  assign nG_101_38 = nG_101_70 | (nP_101_70 & nG_69_38);
  assign nP_101_38 = nP_101_70 & nP_69_38;
  assign nG_100_37 = nG_100_69 | (nP_100_69 & nG_68_37);
  assign nP_100_37 = nP_100_69 & nP_68_37;
  assign nG_99_36 = nG_99_68 | (nP_99_68 & nG_67_36);
  assign nP_99_36 = nP_99_68 & nP_67_36;
  assign nG_98_35 = nG_98_67 | (nP_98_67 & nG_66_35);
  assign nP_98_35 = nP_98_67 & nP_66_35;
  assign nG_97_34 = nG_97_66 | (nP_97_66 & nG_65_34);
  assign nP_97_34 = nP_97_66 & nP_65_34;
  assign nG_96_33 = nG_96_65 | (nP_96_65 & nG_64_33);
  assign nP_96_33 = nP_96_65 & nP_64_33;
  assign nG_95_32 = nG_95_64 | (nP_95_64 & nG_63_32);
  assign nP_95_32 = nP_95_64 & nP_63_32;
  assign nG_94_31 = nG_94_63 | (nP_94_63 & nG_62_31);
  assign nP_94_31 = nP_94_63 & nP_62_31;
  assign nG_93_30 = nG_93_62 | (nP_93_62 & nG_61_30);
  assign nP_93_30 = nP_93_62 & nP_61_30;
  assign nG_92_29 = nG_92_61 | (nP_92_61 & nG_60_29);
  assign nP_92_29 = nP_92_61 & nP_60_29;
  assign nG_91_28 = nG_91_60 | (nP_91_60 & nG_59_28);
  assign nP_91_28 = nP_91_60 & nP_59_28;
  assign nG_90_27 = nG_90_59 | (nP_90_59 & nG_58_27);
  assign nP_90_27 = nP_90_59 & nP_58_27;
  assign nG_89_26 = nG_89_58 | (nP_89_58 & nG_57_26);
  assign nP_89_26 = nP_89_58 & nP_57_26;
  assign nG_88_25 = nG_88_57 | (nP_88_57 & nG_56_25);
  assign nP_88_25 = nP_88_57 & nP_56_25;
  assign nG_87_24 = nG_87_56 | (nP_87_56 & nG_55_24);
  assign nP_87_24 = nP_87_56 & nP_55_24;
  assign nG_86_23 = nG_86_55 | (nP_86_55 & nG_54_23);
  assign nP_86_23 = nP_86_55 & nP_54_23;
  assign nG_85_22 = nG_85_54 | (nP_85_54 & nG_53_22);
  assign nP_85_22 = nP_85_54 & nP_53_22;
  assign nG_84_21 = nG_84_53 | (nP_84_53 & nG_52_21);
  assign nP_84_21 = nP_84_53 & nP_52_21;
  assign nG_83_20 = nG_83_52 | (nP_83_52 & nG_51_20);
  assign nP_83_20 = nP_83_52 & nP_51_20;
  assign nG_82_19 = nG_82_51 | (nP_82_51 & nG_50_19);
  assign nP_82_19 = nP_82_51 & nP_50_19;
  assign nG_81_18 = nG_81_50 | (nP_81_50 & nG_49_18);
  assign nP_81_18 = nP_81_50 & nP_49_18;
  assign nG_80_17 = nG_80_49 | (nP_80_49 & nG_48_17);
  assign nP_80_17 = nP_80_49 & nP_48_17;
  assign nG_79_16 = nG_79_48 | (nP_79_48 & nG_47_16);
  assign nP_79_16 = nP_79_48 & nP_47_16;
  assign nG_78_15 = nG_78_47 | (nP_78_47 & nG_46_15);
  assign nP_78_15 = nP_78_47 & nP_46_15;
  assign nG_77_14 = nG_77_46 | (nP_77_46 & nG_45_14);
  assign nP_77_14 = nP_77_46 & nP_45_14;
  assign nG_76_13 = nG_76_45 | (nP_76_45 & nG_44_13);
  assign nP_76_13 = nP_76_45 & nP_44_13;
  assign nG_75_12 = nG_75_44 | (nP_75_44 & nG_43_12);
  assign nP_75_12 = nP_75_44 & nP_43_12;
  assign nG_74_11 = nG_74_43 | (nP_74_43 & nG_42_11);
  assign nP_74_11 = nP_74_43 & nP_42_11;
  assign nG_73_10 = nG_73_42 | (nP_73_42 & nG_41_10);
  assign nP_73_10 = nP_73_42 & nP_41_10;
  assign nG_72_9 = nG_72_41 | (nP_72_41 & nG_40_9);
  assign nP_72_9 = nP_72_41 & nP_40_9;
  assign nG_71_8 = nG_71_40 | (nP_71_40 & nG_39_8);
  assign nP_71_8 = nP_71_40 & nP_39_8;
  assign nG_70_7 = nG_70_39 | (nP_70_39 & nG_38_7);
  assign nP_70_7 = nP_70_39 & nP_38_7;
  assign nG_69_6 = nG_69_38 | (nP_69_38 & nG_37_6);
  assign nP_69_6 = nP_69_38 & nP_37_6;
  assign nG_68_5 = nG_68_37 | (nP_68_37 & nG_36_5);
  assign nP_68_5 = nP_68_37 & nP_36_5;
  assign nG_67_4 = nG_67_36 | (nP_67_36 & nG_35_4);
  assign nP_67_4 = nP_67_36 & nP_35_4;
  assign nG_66_3 = nG_66_35 | (nP_66_35 & nG_34_3);
  assign nP_66_3 = nP_66_35 & nP_34_3;
  assign nG_65_2 = nG_65_34 | (nP_65_34 & nG_33_2);
  assign nP_65_2 = nP_65_34 & nP_33_2;
  assign nG_64_1 = nG_64_33 | (nP_64_33 & nG_32_1);
  assign nP_64_1 = nP_64_33 & nP_32_1;
  assign nG_63_0 = nG_63_32 | (nP_63_32 & nG_31_0);
  assign nP_63_0 = nP_63_32 & nP_31_0;
  assign nG_62_0 = nG_62_31 | (nP_62_31 & nG_30_0);
  assign nP_62_0 = nP_62_31 & nP_30_0;
  assign nG_61_0 = nG_61_30 | (nP_61_30 & nG_29_0);
  assign nP_61_0 = nP_61_30 & nP_29_0;
  assign nG_60_0 = nG_60_29 | (nP_60_29 & nG_28_0);
  assign nP_60_0 = nP_60_29 & nP_28_0;
  assign nG_59_0 = nG_59_28 | (nP_59_28 & nG_27_0);
  assign nP_59_0 = nP_59_28 & nP_27_0;
  assign nG_58_0 = nG_58_27 | (nP_58_27 & nG_26_0);
  assign nP_58_0 = nP_58_27 & nP_26_0;
  assign nG_57_0 = nG_57_26 | (nP_57_26 & nG_25_0);
  assign nP_57_0 = nP_57_26 & nP_25_0;
  assign nG_56_0 = nG_56_25 | (nP_56_25 & nG_24_0);
  assign nP_56_0 = nP_56_25 & nP_24_0;
  assign nG_55_0 = nG_55_24 | (nP_55_24 & nG_23_0);
  assign nP_55_0 = nP_55_24 & nP_23_0;
  assign nG_54_0 = nG_54_23 | (nP_54_23 & nG_22_0);
  assign nP_54_0 = nP_54_23 & nP_22_0;
  assign nG_53_0 = nG_53_22 | (nP_53_22 & nG_21_0);
  assign nP_53_0 = nP_53_22 & nP_21_0;
  assign nG_52_0 = nG_52_21 | (nP_52_21 & nG_20_0);
  assign nP_52_0 = nP_52_21 & nP_20_0;
  assign nG_51_0 = nG_51_20 | (nP_51_20 & nG_19_0);
  assign nP_51_0 = nP_51_20 & nP_19_0;
  assign nG_50_0 = nG_50_19 | (nP_50_19 & nG_18_0);
  assign nP_50_0 = nP_50_19 & nP_18_0;
  assign nG_49_0 = nG_49_18 | (nP_49_18 & nG_17_0);
  assign nP_49_0 = nP_49_18 & nP_17_0;
  assign nG_48_0 = nG_48_17 | (nP_48_17 & nG_16_0);
  assign nP_48_0 = nP_48_17 & nP_16_0;
  assign nG_47_0 = nG_47_16 | (nP_47_16 & nG_15_0);
  assign nP_47_0 = nP_47_16 & nP_15_0;
  assign nG_46_0 = nG_46_15 | (nP_46_15 & nG_14_0);
  assign nP_46_0 = nP_46_15 & nP_14_0;
  assign nG_45_0 = nG_45_14 | (nP_45_14 & nG_13_0);
  assign nP_45_0 = nP_45_14 & nP_13_0;
  assign nG_44_0 = nG_44_13 | (nP_44_13 & nG_12_0);
  assign nP_44_0 = nP_44_13 & nP_12_0;
  assign nG_43_0 = nG_43_12 | (nP_43_12 & nG_11_0);
  assign nP_43_0 = nP_43_12 & nP_11_0;
  assign nG_42_0 = nG_42_11 | (nP_42_11 & nG_10_0);
  assign nP_42_0 = nP_42_11 & nP_10_0;
  assign nG_41_0 = nG_41_10 | (nP_41_10 & nG_9_0);
  assign nP_41_0 = nP_41_10 & nP_9_0;
  assign nG_40_0 = nG_40_9 | (nP_40_9 & nG_8_0);
  assign nP_40_0 = nP_40_9 & nP_8_0;
  assign nG_39_0 = nG_39_8 | (nP_39_8 & nG_7_0);
  assign nP_39_0 = nP_39_8 & nP_7_0;
  assign nG_38_0 = nG_38_7 | (nP_38_7 & nG_6_0);
  assign nP_38_0 = nP_38_7 & nP_6_0;
  assign nG_37_0 = nG_37_6 | (nP_37_6 & nG_5_0);
  assign nP_37_0 = nP_37_6 & nP_5_0;
  assign nG_36_0 = nG_36_5 | (nP_36_5 & nG_4_0);
  assign nP_36_0 = nP_36_5 & nP_4_0;
  assign nG_35_0 = nG_35_4 | (nP_35_4 & nG_3_0);
  assign nP_35_0 = nP_35_4 & nP_3_0;
  assign nG_34_0 = nG_34_3 | (nP_34_3 & nG_2_0);
  assign nP_34_0 = nP_34_3 & nP_2_0;
  assign nG_33_0 = nG_33_2 | (nP_33_2 & nG_1_0);
  assign nP_33_0 = nP_33_2 & nP_1_0;
  assign nG_32_0 = nG_32_1 | (nP_32_1 & nG_0_0);
  assign nP_32_0 = nP_32_1 & nP_0_0;

  assign nG_127_0 = nG_127_64 | (nP_127_64 & nG_63_0);
  assign nP_127_0 = nP_127_64 & nP_63_0;
  assign nG_126_0 = nG_126_63 | (nP_126_63 & nG_62_0);
  assign nP_126_0 = nP_126_63 & nP_62_0;
  assign nG_125_0 = nG_125_62 | (nP_125_62 & nG_61_0);
  assign nP_125_0 = nP_125_62 & nP_61_0;
  assign nG_124_0 = nG_124_61 | (nP_124_61 & nG_60_0);
  assign nP_124_0 = nP_124_61 & nP_60_0;
  assign nG_123_0 = nG_123_60 | (nP_123_60 & nG_59_0);
  assign nP_123_0 = nP_123_60 & nP_59_0;
  assign nG_122_0 = nG_122_59 | (nP_122_59 & nG_58_0);
  assign nP_122_0 = nP_122_59 & nP_58_0;
  assign nG_121_0 = nG_121_58 | (nP_121_58 & nG_57_0);
  assign nP_121_0 = nP_121_58 & nP_57_0;
  assign nG_120_0 = nG_120_57 | (nP_120_57 & nG_56_0);
  assign nP_120_0 = nP_120_57 & nP_56_0;
  assign nG_119_0 = nG_119_56 | (nP_119_56 & nG_55_0);
  assign nP_119_0 = nP_119_56 & nP_55_0;
  assign nG_118_0 = nG_118_55 | (nP_118_55 & nG_54_0);
  assign nP_118_0 = nP_118_55 & nP_54_0;
  assign nG_117_0 = nG_117_54 | (nP_117_54 & nG_53_0);
  assign nP_117_0 = nP_117_54 & nP_53_0;
  assign nG_116_0 = nG_116_53 | (nP_116_53 & nG_52_0);
  assign nP_116_0 = nP_116_53 & nP_52_0;
  assign nG_115_0 = nG_115_52 | (nP_115_52 & nG_51_0);
  assign nP_115_0 = nP_115_52 & nP_51_0;
  assign nG_114_0 = nG_114_51 | (nP_114_51 & nG_50_0);
  assign nP_114_0 = nP_114_51 & nP_50_0;
  assign nG_113_0 = nG_113_50 | (nP_113_50 & nG_49_0);
  assign nP_113_0 = nP_113_50 & nP_49_0;
  assign nG_112_0 = nG_112_49 | (nP_112_49 & nG_48_0);
  assign nP_112_0 = nP_112_49 & nP_48_0;
  assign nG_111_0 = nG_111_48 | (nP_111_48 & nG_47_0);
  assign nP_111_0 = nP_111_48 & nP_47_0;
  assign nG_110_0 = nG_110_47 | (nP_110_47 & nG_46_0);
  assign nP_110_0 = nP_110_47 & nP_46_0;
  assign nG_109_0 = nG_109_46 | (nP_109_46 & nG_45_0);
  assign nP_109_0 = nP_109_46 & nP_45_0;
  assign nG_108_0 = nG_108_45 | (nP_108_45 & nG_44_0);
  assign nP_108_0 = nP_108_45 & nP_44_0;
  assign nG_107_0 = nG_107_44 | (nP_107_44 & nG_43_0);
  assign nP_107_0 = nP_107_44 & nP_43_0;
  assign nG_106_0 = nG_106_43 | (nP_106_43 & nG_42_0);
  assign nP_106_0 = nP_106_43 & nP_42_0;
  assign nG_105_0 = nG_105_42 | (nP_105_42 & nG_41_0);
  assign nP_105_0 = nP_105_42 & nP_41_0;
  assign nG_104_0 = nG_104_41 | (nP_104_41 & nG_40_0);
  assign nP_104_0 = nP_104_41 & nP_40_0;
  assign nG_103_0 = nG_103_40 | (nP_103_40 & nG_39_0);
  assign nP_103_0 = nP_103_40 & nP_39_0;
  assign nG_102_0 = nG_102_39 | (nP_102_39 & nG_38_0);
  assign nP_102_0 = nP_102_39 & nP_38_0;
  assign nG_101_0 = nG_101_38 | (nP_101_38 & nG_37_0);
  assign nP_101_0 = nP_101_38 & nP_37_0;
  assign nG_100_0 = nG_100_37 | (nP_100_37 & nG_36_0);
  assign nP_100_0 = nP_100_37 & nP_36_0;
  assign nG_99_0 = nG_99_36 | (nP_99_36 & nG_35_0);
  assign nP_99_0 = nP_99_36 & nP_35_0;
  assign nG_98_0 = nG_98_35 | (nP_98_35 & nG_34_0);
  assign nP_98_0 = nP_98_35 & nP_34_0;
  assign nG_97_0 = nG_97_34 | (nP_97_34 & nG_33_0);
  assign nP_97_0 = nP_97_34 & nP_33_0;
  assign nG_96_0 = nG_96_33 | (nP_96_33 & nG_32_0);
  assign nP_96_0 = nP_96_33 & nP_32_0;
  assign nG_95_0 = nG_95_32 | (nP_95_32 & nG_31_0);
  assign nP_95_0 = nP_95_32 & nP_31_0;
  assign nG_94_0 = nG_94_31 | (nP_94_31 & nG_30_0);
  assign nP_94_0 = nP_94_31 & nP_30_0;
  assign nG_93_0 = nG_93_30 | (nP_93_30 & nG_29_0);
  assign nP_93_0 = nP_93_30 & nP_29_0;
  assign nG_92_0 = nG_92_29 | (nP_92_29 & nG_28_0);
  assign nP_92_0 = nP_92_29 & nP_28_0;
  assign nG_91_0 = nG_91_28 | (nP_91_28 & nG_27_0);
  assign nP_91_0 = nP_91_28 & nP_27_0;
  assign nG_90_0 = nG_90_27 | (nP_90_27 & nG_26_0);
  assign nP_90_0 = nP_90_27 & nP_26_0;
  assign nG_89_0 = nG_89_26 | (nP_89_26 & nG_25_0);
  assign nP_89_0 = nP_89_26 & nP_25_0;
  assign nG_88_0 = nG_88_25 | (nP_88_25 & nG_24_0);
  assign nP_88_0 = nP_88_25 & nP_24_0;
  assign nG_87_0 = nG_87_24 | (nP_87_24 & nG_23_0);
  assign nP_87_0 = nP_87_24 & nP_23_0;
  assign nG_86_0 = nG_86_23 | (nP_86_23 & nG_22_0);
  assign nP_86_0 = nP_86_23 & nP_22_0;
  assign nG_85_0 = nG_85_22 | (nP_85_22 & nG_21_0);
  assign nP_85_0 = nP_85_22 & nP_21_0;
  assign nG_84_0 = nG_84_21 | (nP_84_21 & nG_20_0);
  assign nP_84_0 = nP_84_21 & nP_20_0;
  assign nG_83_0 = nG_83_20 | (nP_83_20 & nG_19_0);
  assign nP_83_0 = nP_83_20 & nP_19_0;
  assign nG_82_0 = nG_82_19 | (nP_82_19 & nG_18_0);
  assign nP_82_0 = nP_82_19 & nP_18_0;
  assign nG_81_0 = nG_81_18 | (nP_81_18 & nG_17_0);
  assign nP_81_0 = nP_81_18 & nP_17_0;
  assign nG_80_0 = nG_80_17 | (nP_80_17 & nG_16_0);
  assign nP_80_0 = nP_80_17 & nP_16_0;
  assign nG_79_0 = nG_79_16 | (nP_79_16 & nG_15_0);
  assign nP_79_0 = nP_79_16 & nP_15_0;
  assign nG_78_0 = nG_78_15 | (nP_78_15 & nG_14_0);
  assign nP_78_0 = nP_78_15 & nP_14_0;
  assign nG_77_0 = nG_77_14 | (nP_77_14 & nG_13_0);
  assign nP_77_0 = nP_77_14 & nP_13_0;
  assign nG_76_0 = nG_76_13 | (nP_76_13 & nG_12_0);
  assign nP_76_0 = nP_76_13 & nP_12_0;
  assign nG_75_0 = nG_75_12 | (nP_75_12 & nG_11_0);
  assign nP_75_0 = nP_75_12 & nP_11_0;
  assign nG_74_0 = nG_74_11 | (nP_74_11 & nG_10_0);
  assign nP_74_0 = nP_74_11 & nP_10_0;
  assign nG_73_0 = nG_73_10 | (nP_73_10 & nG_9_0);
  assign nP_73_0 = nP_73_10 & nP_9_0;
  assign nG_72_0 = nG_72_9 | (nP_72_9 & nG_8_0);
  assign nP_72_0 = nP_72_9 & nP_8_0;
  assign nG_71_0 = nG_71_8 | (nP_71_8 & nG_7_0);
  assign nP_71_0 = nP_71_8 & nP_7_0;
  assign nG_70_0 = nG_70_7 | (nP_70_7 & nG_6_0);
  assign nP_70_0 = nP_70_7 & nP_6_0;
  assign nG_69_0 = nG_69_6 | (nP_69_6 & nG_5_0);
  assign nP_69_0 = nP_69_6 & nP_5_0;
  assign nG_68_0 = nG_68_5 | (nP_68_5 & nG_4_0);
  assign nP_68_0 = nP_68_5 & nP_4_0;
  assign nG_67_0 = nG_67_4 | (nP_67_4 & nG_3_0);
  assign nP_67_0 = nP_67_4 & nP_3_0;
  assign nG_66_0 = nG_66_3 | (nP_66_3 & nG_2_0);
  assign nP_66_0 = nP_66_3 & nP_2_0;
  assign nG_65_0 = nG_65_2 | (nP_65_2 & nG_1_0);
  assign nP_65_0 = nP_65_2 & nP_1_0;
  assign nG_64_0 = nG_64_1 | (nP_64_1 & nG_0_0);
  assign nP_64_0 = nP_64_1 & nP_0_0;

  assign nC_0 = in_CI;
  assign nC_1 = nG_0_0 | (nP_0_0 & in_CI);
  assign nC_2 = nG_1_0 | (nP_1_0 & in_CI);
  assign nC_3 = nG_2_0 | (nP_2_0 & in_CI);
  assign nC_4 = nG_3_0 | (nP_3_0 & in_CI);
  assign nC_5 = nG_4_0 | (nP_4_0 & in_CI);
  assign nC_6 = nG_5_0 | (nP_5_0 & in_CI);
  assign nC_7 = nG_6_0 | (nP_6_0 & in_CI);
  assign nC_8 = nG_7_0 | (nP_7_0 & in_CI);
  assign nC_9 = nG_8_0 | (nP_8_0 & in_CI);
  assign nC_10 = nG_9_0 | (nP_9_0 & in_CI);
  assign nC_11 = nG_10_0 | (nP_10_0 & in_CI);
  assign nC_12 = nG_11_0 | (nP_11_0 & in_CI);
  assign nC_13 = nG_12_0 | (nP_12_0 & in_CI);
  assign nC_14 = nG_13_0 | (nP_13_0 & in_CI);
  assign nC_15 = nG_14_0 | (nP_14_0 & in_CI);
  assign nC_16 = nG_15_0 | (nP_15_0 & in_CI);
  assign nC_17 = nG_16_0 | (nP_16_0 & in_CI);
  assign nC_18 = nG_17_0 | (nP_17_0 & in_CI);
  assign nC_19 = nG_18_0 | (nP_18_0 & in_CI);
  assign nC_20 = nG_19_0 | (nP_19_0 & in_CI);
  assign nC_21 = nG_20_0 | (nP_20_0 & in_CI);
  assign nC_22 = nG_21_0 | (nP_21_0 & in_CI);
  assign nC_23 = nG_22_0 | (nP_22_0 & in_CI);
  assign nC_24 = nG_23_0 | (nP_23_0 & in_CI);
  assign nC_25 = nG_24_0 | (nP_24_0 & in_CI);
  assign nC_26 = nG_25_0 | (nP_25_0 & in_CI);
  assign nC_27 = nG_26_0 | (nP_26_0 & in_CI);
  assign nC_28 = nG_27_0 | (nP_27_0 & in_CI);
  assign nC_29 = nG_28_0 | (nP_28_0 & in_CI);
  assign nC_30 = nG_29_0 | (nP_29_0 & in_CI);
  assign nC_31 = nG_30_0 | (nP_30_0 & in_CI);
  assign nC_32 = nG_31_0 | (nP_31_0 & in_CI);
  assign nC_33 = nG_32_0 | (nP_32_0 & in_CI);
  assign nC_34 = nG_33_0 | (nP_33_0 & in_CI);
  assign nC_35 = nG_34_0 | (nP_34_0 & in_CI);
  assign nC_36 = nG_35_0 | (nP_35_0 & in_CI);
  assign nC_37 = nG_36_0 | (nP_36_0 & in_CI);
  assign nC_38 = nG_37_0 | (nP_37_0 & in_CI);
  assign nC_39 = nG_38_0 | (nP_38_0 & in_CI);
  assign nC_40 = nG_39_0 | (nP_39_0 & in_CI);
  assign nC_41 = nG_40_0 | (nP_40_0 & in_CI);
  assign nC_42 = nG_41_0 | (nP_41_0 & in_CI);
  assign nC_43 = nG_42_0 | (nP_42_0 & in_CI);
  assign nC_44 = nG_43_0 | (nP_43_0 & in_CI);
  assign nC_45 = nG_44_0 | (nP_44_0 & in_CI);
  assign nC_46 = nG_45_0 | (nP_45_0 & in_CI);
  assign nC_47 = nG_46_0 | (nP_46_0 & in_CI);
  assign nC_48 = nG_47_0 | (nP_47_0 & in_CI);
  assign nC_49 = nG_48_0 | (nP_48_0 & in_CI);
  assign nC_50 = nG_49_0 | (nP_49_0 & in_CI);
  assign nC_51 = nG_50_0 | (nP_50_0 & in_CI);
  assign nC_52 = nG_51_0 | (nP_51_0 & in_CI);
  assign nC_53 = nG_52_0 | (nP_52_0 & in_CI);
  assign nC_54 = nG_53_0 | (nP_53_0 & in_CI);
  assign nC_55 = nG_54_0 | (nP_54_0 & in_CI);
  assign nC_56 = nG_55_0 | (nP_55_0 & in_CI);
  assign nC_57 = nG_56_0 | (nP_56_0 & in_CI);
  assign nC_58 = nG_57_0 | (nP_57_0 & in_CI);
  assign nC_59 = nG_58_0 | (nP_58_0 & in_CI);
  assign nC_60 = nG_59_0 | (nP_59_0 & in_CI);
  assign nC_61 = nG_60_0 | (nP_60_0 & in_CI);
  assign nC_62 = nG_61_0 | (nP_61_0 & in_CI);
  assign nC_63 = nG_62_0 | (nP_62_0 & in_CI);
  assign nC_64 = nG_63_0 | (nP_63_0 & in_CI);
  assign nC_65 = nG_64_0 | (nP_64_0 & in_CI);
  assign nC_66 = nG_65_0 | (nP_65_0 & in_CI);
  assign nC_67 = nG_66_0 | (nP_66_0 & in_CI);
  assign nC_68 = nG_67_0 | (nP_67_0 & in_CI);
  assign nC_69 = nG_68_0 | (nP_68_0 & in_CI);
  assign nC_70 = nG_69_0 | (nP_69_0 & in_CI);
  assign nC_71 = nG_70_0 | (nP_70_0 & in_CI);
  assign nC_72 = nG_71_0 | (nP_71_0 & in_CI);
  assign nC_73 = nG_72_0 | (nP_72_0 & in_CI);
  assign nC_74 = nG_73_0 | (nP_73_0 & in_CI);
  assign nC_75 = nG_74_0 | (nP_74_0 & in_CI);
  assign nC_76 = nG_75_0 | (nP_75_0 & in_CI);
  assign nC_77 = nG_76_0 | (nP_76_0 & in_CI);
  assign nC_78 = nG_77_0 | (nP_77_0 & in_CI);
  assign nC_79 = nG_78_0 | (nP_78_0 & in_CI);
  assign nC_80 = nG_79_0 | (nP_79_0 & in_CI);
  assign nC_81 = nG_80_0 | (nP_80_0 & in_CI);
  assign nC_82 = nG_81_0 | (nP_81_0 & in_CI);
  assign nC_83 = nG_82_0 | (nP_82_0 & in_CI);
  assign nC_84 = nG_83_0 | (nP_83_0 & in_CI);
  assign nC_85 = nG_84_0 | (nP_84_0 & in_CI);
  assign nC_86 = nG_85_0 | (nP_85_0 & in_CI);
  assign nC_87 = nG_86_0 | (nP_86_0 & in_CI);
  assign nC_88 = nG_87_0 | (nP_87_0 & in_CI);
  assign nC_89 = nG_88_0 | (nP_88_0 & in_CI);
  assign nC_90 = nG_89_0 | (nP_89_0 & in_CI);
  assign nC_91 = nG_90_0 | (nP_90_0 & in_CI);
  assign nC_92 = nG_91_0 | (nP_91_0 & in_CI);
  assign nC_93 = nG_92_0 | (nP_92_0 & in_CI);
  assign nC_94 = nG_93_0 | (nP_93_0 & in_CI);
  assign nC_95 = nG_94_0 | (nP_94_0 & in_CI);
  assign nC_96 = nG_95_0 | (nP_95_0 & in_CI);
  assign nC_97 = nG_96_0 | (nP_96_0 & in_CI);
  assign nC_98 = nG_97_0 | (nP_97_0 & in_CI);
  assign nC_99 = nG_98_0 | (nP_98_0 & in_CI);
  assign nC_100 = nG_99_0 | (nP_99_0 & in_CI);
  assign nC_101 = nG_100_0 | (nP_100_0 & in_CI);
  assign nC_102 = nG_101_0 | (nP_101_0 & in_CI);
  assign nC_103 = nG_102_0 | (nP_102_0 & in_CI);
  assign nC_104 = nG_103_0 | (nP_103_0 & in_CI);
  assign nC_105 = nG_104_0 | (nP_104_0 & in_CI);
  assign nC_106 = nG_105_0 | (nP_105_0 & in_CI);
  assign nC_107 = nG_106_0 | (nP_106_0 & in_CI);
  assign nC_108 = nG_107_0 | (nP_107_0 & in_CI);
  assign nC_109 = nG_108_0 | (nP_108_0 & in_CI);
  assign nC_110 = nG_109_0 | (nP_109_0 & in_CI);
  assign nC_111 = nG_110_0 | (nP_110_0 & in_CI);
  assign nC_112 = nG_111_0 | (nP_111_0 & in_CI);
  assign nC_113 = nG_112_0 | (nP_112_0 & in_CI);
  assign nC_114 = nG_113_0 | (nP_113_0 & in_CI);
  assign nC_115 = nG_114_0 | (nP_114_0 & in_CI);
  assign nC_116 = nG_115_0 | (nP_115_0 & in_CI);
  assign nC_117 = nG_116_0 | (nP_116_0 & in_CI);
  assign nC_118 = nG_117_0 | (nP_117_0 & in_CI);
  assign nC_119 = nG_118_0 | (nP_118_0 & in_CI);
  assign nC_120 = nG_119_0 | (nP_119_0 & in_CI);
  assign nC_121 = nG_120_0 | (nP_120_0 & in_CI);
  assign nC_122 = nG_121_0 | (nP_121_0 & in_CI);
  assign nC_123 = nG_122_0 | (nP_122_0 & in_CI);
  assign nC_124 = nG_123_0 | (nP_123_0 & in_CI);
  assign nC_125 = nG_124_0 | (nP_124_0 & in_CI);
  assign nC_126 = nG_125_0 | (nP_125_0 & in_CI);
  assign nC_127 = nG_126_0 | (nP_126_0 & in_CI);

  assign out_S[0] = nP_0_0 ^ nC_0;
  assign out_S[1] = nP_1_1 ^ nC_1;
  assign out_S[2] = nP_2_2 ^ nC_2;
  assign out_S[3] = nP_3_3 ^ nC_3;
  assign out_S[4] = nP_4_4 ^ nC_4;
  assign out_S[5] = nP_5_5 ^ nC_5;
  assign out_S[6] = nP_6_6 ^ nC_6;
  assign out_S[7] = nP_7_7 ^ nC_7;
  assign out_S[8] = nP_8_8 ^ nC_8;
  assign out_S[9] = nP_9_9 ^ nC_9;
  assign out_S[10] = nP_10_10 ^ nC_10;
  assign out_S[11] = nP_11_11 ^ nC_11;
  assign out_S[12] = nP_12_12 ^ nC_12;
  assign out_S[13] = nP_13_13 ^ nC_13;
  assign out_S[14] = nP_14_14 ^ nC_14;
  assign out_S[15] = nP_15_15 ^ nC_15;
  assign out_S[16] = nP_16_16 ^ nC_16;
  assign out_S[17] = nP_17_17 ^ nC_17;
  assign out_S[18] = nP_18_18 ^ nC_18;
  assign out_S[19] = nP_19_19 ^ nC_19;
  assign out_S[20] = nP_20_20 ^ nC_20;
  assign out_S[21] = nP_21_21 ^ nC_21;
  assign out_S[22] = nP_22_22 ^ nC_22;
  assign out_S[23] = nP_23_23 ^ nC_23;
  assign out_S[24] = nP_24_24 ^ nC_24;
  assign out_S[25] = nP_25_25 ^ nC_25;
  assign out_S[26] = nP_26_26 ^ nC_26;
  assign out_S[27] = nP_27_27 ^ nC_27;
  assign out_S[28] = nP_28_28 ^ nC_28;
  assign out_S[29] = nP_29_29 ^ nC_29;
  assign out_S[30] = nP_30_30 ^ nC_30;
  assign out_S[31] = nP_31_31 ^ nC_31;
  assign out_S[32] = nP_32_32 ^ nC_32;
  assign out_S[33] = nP_33_33 ^ nC_33;
  assign out_S[34] = nP_34_34 ^ nC_34;
  assign out_S[35] = nP_35_35 ^ nC_35;
  assign out_S[36] = nP_36_36 ^ nC_36;
  assign out_S[37] = nP_37_37 ^ nC_37;
  assign out_S[38] = nP_38_38 ^ nC_38;
  assign out_S[39] = nP_39_39 ^ nC_39;
  assign out_S[40] = nP_40_40 ^ nC_40;
  assign out_S[41] = nP_41_41 ^ nC_41;
  assign out_S[42] = nP_42_42 ^ nC_42;
  assign out_S[43] = nP_43_43 ^ nC_43;
  assign out_S[44] = nP_44_44 ^ nC_44;
  assign out_S[45] = nP_45_45 ^ nC_45;
  assign out_S[46] = nP_46_46 ^ nC_46;
  assign out_S[47] = nP_47_47 ^ nC_47;
  assign out_S[48] = nP_48_48 ^ nC_48;
  assign out_S[49] = nP_49_49 ^ nC_49;
  assign out_S[50] = nP_50_50 ^ nC_50;
  assign out_S[51] = nP_51_51 ^ nC_51;
  assign out_S[52] = nP_52_52 ^ nC_52;
  assign out_S[53] = nP_53_53 ^ nC_53;
  assign out_S[54] = nP_54_54 ^ nC_54;
  assign out_S[55] = nP_55_55 ^ nC_55;
  assign out_S[56] = nP_56_56 ^ nC_56;
  assign out_S[57] = nP_57_57 ^ nC_57;
  assign out_S[58] = nP_58_58 ^ nC_58;
  assign out_S[59] = nP_59_59 ^ nC_59;
  assign out_S[60] = nP_60_60 ^ nC_60;
  assign out_S[61] = nP_61_61 ^ nC_61;
  assign out_S[62] = nP_62_62 ^ nC_62;
  assign out_S[63] = nP_63_63 ^ nC_63;
  assign out_S[64] = nP_64_64 ^ nC_64;
  assign out_S[65] = nP_65_65 ^ nC_65;
  assign out_S[66] = nP_66_66 ^ nC_66;
  assign out_S[67] = nP_67_67 ^ nC_67;
  assign out_S[68] = nP_68_68 ^ nC_68;
  assign out_S[69] = nP_69_69 ^ nC_69;
  assign out_S[70] = nP_70_70 ^ nC_70;
  assign out_S[71] = nP_71_71 ^ nC_71;
  assign out_S[72] = nP_72_72 ^ nC_72;
  assign out_S[73] = nP_73_73 ^ nC_73;
  assign out_S[74] = nP_74_74 ^ nC_74;
  assign out_S[75] = nP_75_75 ^ nC_75;
  assign out_S[76] = nP_76_76 ^ nC_76;
  assign out_S[77] = nP_77_77 ^ nC_77;
  assign out_S[78] = nP_78_78 ^ nC_78;
  assign out_S[79] = nP_79_79 ^ nC_79;
  assign out_S[80] = nP_80_80 ^ nC_80;
  assign out_S[81] = nP_81_81 ^ nC_81;
  assign out_S[82] = nP_82_82 ^ nC_82;
  assign out_S[83] = nP_83_83 ^ nC_83;
  assign out_S[84] = nP_84_84 ^ nC_84;
  assign out_S[85] = nP_85_85 ^ nC_85;
  assign out_S[86] = nP_86_86 ^ nC_86;
  assign out_S[87] = nP_87_87 ^ nC_87;
  assign out_S[88] = nP_88_88 ^ nC_88;
  assign out_S[89] = nP_89_89 ^ nC_89;
  assign out_S[90] = nP_90_90 ^ nC_90;
  assign out_S[91] = nP_91_91 ^ nC_91;
  assign out_S[92] = nP_92_92 ^ nC_92;
  assign out_S[93] = nP_93_93 ^ nC_93;
  assign out_S[94] = nP_94_94 ^ nC_94;
  assign out_S[95] = nP_95_95 ^ nC_95;
  assign out_S[96] = nP_96_96 ^ nC_96;
  assign out_S[97] = nP_97_97 ^ nC_97;
  assign out_S[98] = nP_98_98 ^ nC_98;
  assign out_S[99] = nP_99_99 ^ nC_99;
  assign out_S[100] = nP_100_100 ^ nC_100;
  assign out_S[101] = nP_101_101 ^ nC_101;
  assign out_S[102] = nP_102_102 ^ nC_102;
  assign out_S[103] = nP_103_103 ^ nC_103;
  assign out_S[104] = nP_104_104 ^ nC_104;
  assign out_S[105] = nP_105_105 ^ nC_105;
  assign out_S[106] = nP_106_106 ^ nC_106;
  assign out_S[107] = nP_107_107 ^ nC_107;
  assign out_S[108] = nP_108_108 ^ nC_108;
  assign out_S[109] = nP_109_109 ^ nC_109;
  assign out_S[110] = nP_110_110 ^ nC_110;
  assign out_S[111] = nP_111_111 ^ nC_111;
  assign out_S[112] = nP_112_112 ^ nC_112;
  assign out_S[113] = nP_113_113 ^ nC_113;
  assign out_S[114] = nP_114_114 ^ nC_114;
  assign out_S[115] = nP_115_115 ^ nC_115;
  assign out_S[116] = nP_116_116 ^ nC_116;
  assign out_S[117] = nP_117_117 ^ nC_117;
  assign out_S[118] = nP_118_118 ^ nC_118;
  assign out_S[119] = nP_119_119 ^ nC_119;
  assign out_S[120] = nP_120_120 ^ nC_120;
  assign out_S[121] = nP_121_121 ^ nC_121;
  assign out_S[122] = nP_122_122 ^ nC_122;
  assign out_S[123] = nP_123_123 ^ nC_123;
  assign out_S[124] = nP_124_124 ^ nC_124;
  assign out_S[125] = nP_125_125 ^ nC_125;
  assign out_S[126] = nP_126_126 ^ nC_126;
  assign out_S[127] = nP_127_127 ^ nC_127;
  assign out_CO = nG_127_0 | (nP_127_0 & in_CI);
endmodule

