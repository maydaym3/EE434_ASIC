module VHA (in_A, in_B, out_S, out_CO);
  input in_A, in_B;
  output out_S, out_CO;

  assign out_S = in_A ^ in_B;
  assign out_CO = in_A & in_B;
endmodule

module VFA (in_A, in_B, in_CI, out_S, out_CO);
  input in_A, in_B, in_CI;
  output out_S, out_CO;

  assign out_S = in_A ^ in_B ^ in_CI;
  assign out_CO = (in_A & in_B) | (in_B & in_CI) | (in_CI & in_A);
endmodule



module VCondSumAdder_256 (in_A, in_B, in_CI, out_S, out_CO);
  input [255:0] in_A, in_B;
  input in_CI;
  output [255:0] out_S;
  output out_CO;

  VHA U_st1_b0_c0 (.in_A(in_A[0]), .in_B(in_B[0]), .out_S(nS_st1_b0_c0), .out_CO(nC_st1_b0_c0));
  VFA U_st1_b0_c1 (.in_A(in_A[0]), .in_B(in_B[0]), .in_CI(1'b1), .out_S(nS_st1_b0_c1), .out_CO(nC_st1_b0_c1));
  VHA U_st1_b1_c0 (.in_A(in_A[1]), .in_B(in_B[1]), .out_S(nS_st1_b1_c0), .out_CO(nC_st1_b1_c0));
  VFA U_st1_b1_c1 (.in_A(in_A[1]), .in_B(in_B[1]), .in_CI(1'b1), .out_S(nS_st1_b1_c1), .out_CO(nC_st1_b1_c1));
  VHA U_st1_b2_c0 (.in_A(in_A[2]), .in_B(in_B[2]), .out_S(nS_st1_b2_c0), .out_CO(nC_st1_b2_c0));
  VFA U_st1_b2_c1 (.in_A(in_A[2]), .in_B(in_B[2]), .in_CI(1'b1), .out_S(nS_st1_b2_c1), .out_CO(nC_st1_b2_c1));
  VHA U_st1_b3_c0 (.in_A(in_A[3]), .in_B(in_B[3]), .out_S(nS_st1_b3_c0), .out_CO(nC_st1_b3_c0));
  VFA U_st1_b3_c1 (.in_A(in_A[3]), .in_B(in_B[3]), .in_CI(1'b1), .out_S(nS_st1_b3_c1), .out_CO(nC_st1_b3_c1));
  VHA U_st1_b4_c0 (.in_A(in_A[4]), .in_B(in_B[4]), .out_S(nS_st1_b4_c0), .out_CO(nC_st1_b4_c0));
  VFA U_st1_b4_c1 (.in_A(in_A[4]), .in_B(in_B[4]), .in_CI(1'b1), .out_S(nS_st1_b4_c1), .out_CO(nC_st1_b4_c1));
  VHA U_st1_b5_c0 (.in_A(in_A[5]), .in_B(in_B[5]), .out_S(nS_st1_b5_c0), .out_CO(nC_st1_b5_c0));
  VFA U_st1_b5_c1 (.in_A(in_A[5]), .in_B(in_B[5]), .in_CI(1'b1), .out_S(nS_st1_b5_c1), .out_CO(nC_st1_b5_c1));
  VHA U_st1_b6_c0 (.in_A(in_A[6]), .in_B(in_B[6]), .out_S(nS_st1_b6_c0), .out_CO(nC_st1_b6_c0));
  VFA U_st1_b6_c1 (.in_A(in_A[6]), .in_B(in_B[6]), .in_CI(1'b1), .out_S(nS_st1_b6_c1), .out_CO(nC_st1_b6_c1));
  VHA U_st1_b7_c0 (.in_A(in_A[7]), .in_B(in_B[7]), .out_S(nS_st1_b7_c0), .out_CO(nC_st1_b7_c0));
  VFA U_st1_b7_c1 (.in_A(in_A[7]), .in_B(in_B[7]), .in_CI(1'b1), .out_S(nS_st1_b7_c1), .out_CO(nC_st1_b7_c1));
  VHA U_st1_b8_c0 (.in_A(in_A[8]), .in_B(in_B[8]), .out_S(nS_st1_b8_c0), .out_CO(nC_st1_b8_c0));
  VFA U_st1_b8_c1 (.in_A(in_A[8]), .in_B(in_B[8]), .in_CI(1'b1), .out_S(nS_st1_b8_c1), .out_CO(nC_st1_b8_c1));
  VHA U_st1_b9_c0 (.in_A(in_A[9]), .in_B(in_B[9]), .out_S(nS_st1_b9_c0), .out_CO(nC_st1_b9_c0));
  VFA U_st1_b9_c1 (.in_A(in_A[9]), .in_B(in_B[9]), .in_CI(1'b1), .out_S(nS_st1_b9_c1), .out_CO(nC_st1_b9_c1));
  VHA U_st1_b10_c0 (.in_A(in_A[10]), .in_B(in_B[10]), .out_S(nS_st1_b10_c0), .out_CO(nC_st1_b10_c0));
  VFA U_st1_b10_c1 (.in_A(in_A[10]), .in_B(in_B[10]), .in_CI(1'b1), .out_S(nS_st1_b10_c1), .out_CO(nC_st1_b10_c1));
  VHA U_st1_b11_c0 (.in_A(in_A[11]), .in_B(in_B[11]), .out_S(nS_st1_b11_c0), .out_CO(nC_st1_b11_c0));
  VFA U_st1_b11_c1 (.in_A(in_A[11]), .in_B(in_B[11]), .in_CI(1'b1), .out_S(nS_st1_b11_c1), .out_CO(nC_st1_b11_c1));
  VHA U_st1_b12_c0 (.in_A(in_A[12]), .in_B(in_B[12]), .out_S(nS_st1_b12_c0), .out_CO(nC_st1_b12_c0));
  VFA U_st1_b12_c1 (.in_A(in_A[12]), .in_B(in_B[12]), .in_CI(1'b1), .out_S(nS_st1_b12_c1), .out_CO(nC_st1_b12_c1));
  VHA U_st1_b13_c0 (.in_A(in_A[13]), .in_B(in_B[13]), .out_S(nS_st1_b13_c0), .out_CO(nC_st1_b13_c0));
  VFA U_st1_b13_c1 (.in_A(in_A[13]), .in_B(in_B[13]), .in_CI(1'b1), .out_S(nS_st1_b13_c1), .out_CO(nC_st1_b13_c1));
  VHA U_st1_b14_c0 (.in_A(in_A[14]), .in_B(in_B[14]), .out_S(nS_st1_b14_c0), .out_CO(nC_st1_b14_c0));
  VFA U_st1_b14_c1 (.in_A(in_A[14]), .in_B(in_B[14]), .in_CI(1'b1), .out_S(nS_st1_b14_c1), .out_CO(nC_st1_b14_c1));
  VHA U_st1_b15_c0 (.in_A(in_A[15]), .in_B(in_B[15]), .out_S(nS_st1_b15_c0), .out_CO(nC_st1_b15_c0));
  VFA U_st1_b15_c1 (.in_A(in_A[15]), .in_B(in_B[15]), .in_CI(1'b1), .out_S(nS_st1_b15_c1), .out_CO(nC_st1_b15_c1));
  VHA U_st1_b16_c0 (.in_A(in_A[16]), .in_B(in_B[16]), .out_S(nS_st1_b16_c0), .out_CO(nC_st1_b16_c0));
  VFA U_st1_b16_c1 (.in_A(in_A[16]), .in_B(in_B[16]), .in_CI(1'b1), .out_S(nS_st1_b16_c1), .out_CO(nC_st1_b16_c1));
  VHA U_st1_b17_c0 (.in_A(in_A[17]), .in_B(in_B[17]), .out_S(nS_st1_b17_c0), .out_CO(nC_st1_b17_c0));
  VFA U_st1_b17_c1 (.in_A(in_A[17]), .in_B(in_B[17]), .in_CI(1'b1), .out_S(nS_st1_b17_c1), .out_CO(nC_st1_b17_c1));
  VHA U_st1_b18_c0 (.in_A(in_A[18]), .in_B(in_B[18]), .out_S(nS_st1_b18_c0), .out_CO(nC_st1_b18_c0));
  VFA U_st1_b18_c1 (.in_A(in_A[18]), .in_B(in_B[18]), .in_CI(1'b1), .out_S(nS_st1_b18_c1), .out_CO(nC_st1_b18_c1));
  VHA U_st1_b19_c0 (.in_A(in_A[19]), .in_B(in_B[19]), .out_S(nS_st1_b19_c0), .out_CO(nC_st1_b19_c0));
  VFA U_st1_b19_c1 (.in_A(in_A[19]), .in_B(in_B[19]), .in_CI(1'b1), .out_S(nS_st1_b19_c1), .out_CO(nC_st1_b19_c1));
  VHA U_st1_b20_c0 (.in_A(in_A[20]), .in_B(in_B[20]), .out_S(nS_st1_b20_c0), .out_CO(nC_st1_b20_c0));
  VFA U_st1_b20_c1 (.in_A(in_A[20]), .in_B(in_B[20]), .in_CI(1'b1), .out_S(nS_st1_b20_c1), .out_CO(nC_st1_b20_c1));
  VHA U_st1_b21_c0 (.in_A(in_A[21]), .in_B(in_B[21]), .out_S(nS_st1_b21_c0), .out_CO(nC_st1_b21_c0));
  VFA U_st1_b21_c1 (.in_A(in_A[21]), .in_B(in_B[21]), .in_CI(1'b1), .out_S(nS_st1_b21_c1), .out_CO(nC_st1_b21_c1));
  VHA U_st1_b22_c0 (.in_A(in_A[22]), .in_B(in_B[22]), .out_S(nS_st1_b22_c0), .out_CO(nC_st1_b22_c0));
  VFA U_st1_b22_c1 (.in_A(in_A[22]), .in_B(in_B[22]), .in_CI(1'b1), .out_S(nS_st1_b22_c1), .out_CO(nC_st1_b22_c1));
  VHA U_st1_b23_c0 (.in_A(in_A[23]), .in_B(in_B[23]), .out_S(nS_st1_b23_c0), .out_CO(nC_st1_b23_c0));
  VFA U_st1_b23_c1 (.in_A(in_A[23]), .in_B(in_B[23]), .in_CI(1'b1), .out_S(nS_st1_b23_c1), .out_CO(nC_st1_b23_c1));
  VHA U_st1_b24_c0 (.in_A(in_A[24]), .in_B(in_B[24]), .out_S(nS_st1_b24_c0), .out_CO(nC_st1_b24_c0));
  VFA U_st1_b24_c1 (.in_A(in_A[24]), .in_B(in_B[24]), .in_CI(1'b1), .out_S(nS_st1_b24_c1), .out_CO(nC_st1_b24_c1));
  VHA U_st1_b25_c0 (.in_A(in_A[25]), .in_B(in_B[25]), .out_S(nS_st1_b25_c0), .out_CO(nC_st1_b25_c0));
  VFA U_st1_b25_c1 (.in_A(in_A[25]), .in_B(in_B[25]), .in_CI(1'b1), .out_S(nS_st1_b25_c1), .out_CO(nC_st1_b25_c1));
  VHA U_st1_b26_c0 (.in_A(in_A[26]), .in_B(in_B[26]), .out_S(nS_st1_b26_c0), .out_CO(nC_st1_b26_c0));
  VFA U_st1_b26_c1 (.in_A(in_A[26]), .in_B(in_B[26]), .in_CI(1'b1), .out_S(nS_st1_b26_c1), .out_CO(nC_st1_b26_c1));
  VHA U_st1_b27_c0 (.in_A(in_A[27]), .in_B(in_B[27]), .out_S(nS_st1_b27_c0), .out_CO(nC_st1_b27_c0));
  VFA U_st1_b27_c1 (.in_A(in_A[27]), .in_B(in_B[27]), .in_CI(1'b1), .out_S(nS_st1_b27_c1), .out_CO(nC_st1_b27_c1));
  VHA U_st1_b28_c0 (.in_A(in_A[28]), .in_B(in_B[28]), .out_S(nS_st1_b28_c0), .out_CO(nC_st1_b28_c0));
  VFA U_st1_b28_c1 (.in_A(in_A[28]), .in_B(in_B[28]), .in_CI(1'b1), .out_S(nS_st1_b28_c1), .out_CO(nC_st1_b28_c1));
  VHA U_st1_b29_c0 (.in_A(in_A[29]), .in_B(in_B[29]), .out_S(nS_st1_b29_c0), .out_CO(nC_st1_b29_c0));
  VFA U_st1_b29_c1 (.in_A(in_A[29]), .in_B(in_B[29]), .in_CI(1'b1), .out_S(nS_st1_b29_c1), .out_CO(nC_st1_b29_c1));
  VHA U_st1_b30_c0 (.in_A(in_A[30]), .in_B(in_B[30]), .out_S(nS_st1_b30_c0), .out_CO(nC_st1_b30_c0));
  VFA U_st1_b30_c1 (.in_A(in_A[30]), .in_B(in_B[30]), .in_CI(1'b1), .out_S(nS_st1_b30_c1), .out_CO(nC_st1_b30_c1));
  VHA U_st1_b31_c0 (.in_A(in_A[31]), .in_B(in_B[31]), .out_S(nS_st1_b31_c0), .out_CO(nC_st1_b31_c0));
  VFA U_st1_b31_c1 (.in_A(in_A[31]), .in_B(in_B[31]), .in_CI(1'b1), .out_S(nS_st1_b31_c1), .out_CO(nC_st1_b31_c1));
  VHA U_st1_b32_c0 (.in_A(in_A[32]), .in_B(in_B[32]), .out_S(nS_st1_b32_c0), .out_CO(nC_st1_b32_c0));
  VFA U_st1_b32_c1 (.in_A(in_A[32]), .in_B(in_B[32]), .in_CI(1'b1), .out_S(nS_st1_b32_c1), .out_CO(nC_st1_b32_c1));
  VHA U_st1_b33_c0 (.in_A(in_A[33]), .in_B(in_B[33]), .out_S(nS_st1_b33_c0), .out_CO(nC_st1_b33_c0));
  VFA U_st1_b33_c1 (.in_A(in_A[33]), .in_B(in_B[33]), .in_CI(1'b1), .out_S(nS_st1_b33_c1), .out_CO(nC_st1_b33_c1));
  VHA U_st1_b34_c0 (.in_A(in_A[34]), .in_B(in_B[34]), .out_S(nS_st1_b34_c0), .out_CO(nC_st1_b34_c0));
  VFA U_st1_b34_c1 (.in_A(in_A[34]), .in_B(in_B[34]), .in_CI(1'b1), .out_S(nS_st1_b34_c1), .out_CO(nC_st1_b34_c1));
  VHA U_st1_b35_c0 (.in_A(in_A[35]), .in_B(in_B[35]), .out_S(nS_st1_b35_c0), .out_CO(nC_st1_b35_c0));
  VFA U_st1_b35_c1 (.in_A(in_A[35]), .in_B(in_B[35]), .in_CI(1'b1), .out_S(nS_st1_b35_c1), .out_CO(nC_st1_b35_c1));
  VHA U_st1_b36_c0 (.in_A(in_A[36]), .in_B(in_B[36]), .out_S(nS_st1_b36_c0), .out_CO(nC_st1_b36_c0));
  VFA U_st1_b36_c1 (.in_A(in_A[36]), .in_B(in_B[36]), .in_CI(1'b1), .out_S(nS_st1_b36_c1), .out_CO(nC_st1_b36_c1));
  VHA U_st1_b37_c0 (.in_A(in_A[37]), .in_B(in_B[37]), .out_S(nS_st1_b37_c0), .out_CO(nC_st1_b37_c0));
  VFA U_st1_b37_c1 (.in_A(in_A[37]), .in_B(in_B[37]), .in_CI(1'b1), .out_S(nS_st1_b37_c1), .out_CO(nC_st1_b37_c1));
  VHA U_st1_b38_c0 (.in_A(in_A[38]), .in_B(in_B[38]), .out_S(nS_st1_b38_c0), .out_CO(nC_st1_b38_c0));
  VFA U_st1_b38_c1 (.in_A(in_A[38]), .in_B(in_B[38]), .in_CI(1'b1), .out_S(nS_st1_b38_c1), .out_CO(nC_st1_b38_c1));
  VHA U_st1_b39_c0 (.in_A(in_A[39]), .in_B(in_B[39]), .out_S(nS_st1_b39_c0), .out_CO(nC_st1_b39_c0));
  VFA U_st1_b39_c1 (.in_A(in_A[39]), .in_B(in_B[39]), .in_CI(1'b1), .out_S(nS_st1_b39_c1), .out_CO(nC_st1_b39_c1));
  VHA U_st1_b40_c0 (.in_A(in_A[40]), .in_B(in_B[40]), .out_S(nS_st1_b40_c0), .out_CO(nC_st1_b40_c0));
  VFA U_st1_b40_c1 (.in_A(in_A[40]), .in_B(in_B[40]), .in_CI(1'b1), .out_S(nS_st1_b40_c1), .out_CO(nC_st1_b40_c1));
  VHA U_st1_b41_c0 (.in_A(in_A[41]), .in_B(in_B[41]), .out_S(nS_st1_b41_c0), .out_CO(nC_st1_b41_c0));
  VFA U_st1_b41_c1 (.in_A(in_A[41]), .in_B(in_B[41]), .in_CI(1'b1), .out_S(nS_st1_b41_c1), .out_CO(nC_st1_b41_c1));
  VHA U_st1_b42_c0 (.in_A(in_A[42]), .in_B(in_B[42]), .out_S(nS_st1_b42_c0), .out_CO(nC_st1_b42_c0));
  VFA U_st1_b42_c1 (.in_A(in_A[42]), .in_B(in_B[42]), .in_CI(1'b1), .out_S(nS_st1_b42_c1), .out_CO(nC_st1_b42_c1));
  VHA U_st1_b43_c0 (.in_A(in_A[43]), .in_B(in_B[43]), .out_S(nS_st1_b43_c0), .out_CO(nC_st1_b43_c0));
  VFA U_st1_b43_c1 (.in_A(in_A[43]), .in_B(in_B[43]), .in_CI(1'b1), .out_S(nS_st1_b43_c1), .out_CO(nC_st1_b43_c1));
  VHA U_st1_b44_c0 (.in_A(in_A[44]), .in_B(in_B[44]), .out_S(nS_st1_b44_c0), .out_CO(nC_st1_b44_c0));
  VFA U_st1_b44_c1 (.in_A(in_A[44]), .in_B(in_B[44]), .in_CI(1'b1), .out_S(nS_st1_b44_c1), .out_CO(nC_st1_b44_c1));
  VHA U_st1_b45_c0 (.in_A(in_A[45]), .in_B(in_B[45]), .out_S(nS_st1_b45_c0), .out_CO(nC_st1_b45_c0));
  VFA U_st1_b45_c1 (.in_A(in_A[45]), .in_B(in_B[45]), .in_CI(1'b1), .out_S(nS_st1_b45_c1), .out_CO(nC_st1_b45_c1));
  VHA U_st1_b46_c0 (.in_A(in_A[46]), .in_B(in_B[46]), .out_S(nS_st1_b46_c0), .out_CO(nC_st1_b46_c0));
  VFA U_st1_b46_c1 (.in_A(in_A[46]), .in_B(in_B[46]), .in_CI(1'b1), .out_S(nS_st1_b46_c1), .out_CO(nC_st1_b46_c1));
  VHA U_st1_b47_c0 (.in_A(in_A[47]), .in_B(in_B[47]), .out_S(nS_st1_b47_c0), .out_CO(nC_st1_b47_c0));
  VFA U_st1_b47_c1 (.in_A(in_A[47]), .in_B(in_B[47]), .in_CI(1'b1), .out_S(nS_st1_b47_c1), .out_CO(nC_st1_b47_c1));
  VHA U_st1_b48_c0 (.in_A(in_A[48]), .in_B(in_B[48]), .out_S(nS_st1_b48_c0), .out_CO(nC_st1_b48_c0));
  VFA U_st1_b48_c1 (.in_A(in_A[48]), .in_B(in_B[48]), .in_CI(1'b1), .out_S(nS_st1_b48_c1), .out_CO(nC_st1_b48_c1));
  VHA U_st1_b49_c0 (.in_A(in_A[49]), .in_B(in_B[49]), .out_S(nS_st1_b49_c0), .out_CO(nC_st1_b49_c0));
  VFA U_st1_b49_c1 (.in_A(in_A[49]), .in_B(in_B[49]), .in_CI(1'b1), .out_S(nS_st1_b49_c1), .out_CO(nC_st1_b49_c1));
  VHA U_st1_b50_c0 (.in_A(in_A[50]), .in_B(in_B[50]), .out_S(nS_st1_b50_c0), .out_CO(nC_st1_b50_c0));
  VFA U_st1_b50_c1 (.in_A(in_A[50]), .in_B(in_B[50]), .in_CI(1'b1), .out_S(nS_st1_b50_c1), .out_CO(nC_st1_b50_c1));
  VHA U_st1_b51_c0 (.in_A(in_A[51]), .in_B(in_B[51]), .out_S(nS_st1_b51_c0), .out_CO(nC_st1_b51_c0));
  VFA U_st1_b51_c1 (.in_A(in_A[51]), .in_B(in_B[51]), .in_CI(1'b1), .out_S(nS_st1_b51_c1), .out_CO(nC_st1_b51_c1));
  VHA U_st1_b52_c0 (.in_A(in_A[52]), .in_B(in_B[52]), .out_S(nS_st1_b52_c0), .out_CO(nC_st1_b52_c0));
  VFA U_st1_b52_c1 (.in_A(in_A[52]), .in_B(in_B[52]), .in_CI(1'b1), .out_S(nS_st1_b52_c1), .out_CO(nC_st1_b52_c1));
  VHA U_st1_b53_c0 (.in_A(in_A[53]), .in_B(in_B[53]), .out_S(nS_st1_b53_c0), .out_CO(nC_st1_b53_c0));
  VFA U_st1_b53_c1 (.in_A(in_A[53]), .in_B(in_B[53]), .in_CI(1'b1), .out_S(nS_st1_b53_c1), .out_CO(nC_st1_b53_c1));
  VHA U_st1_b54_c0 (.in_A(in_A[54]), .in_B(in_B[54]), .out_S(nS_st1_b54_c0), .out_CO(nC_st1_b54_c0));
  VFA U_st1_b54_c1 (.in_A(in_A[54]), .in_B(in_B[54]), .in_CI(1'b1), .out_S(nS_st1_b54_c1), .out_CO(nC_st1_b54_c1));
  VHA U_st1_b55_c0 (.in_A(in_A[55]), .in_B(in_B[55]), .out_S(nS_st1_b55_c0), .out_CO(nC_st1_b55_c0));
  VFA U_st1_b55_c1 (.in_A(in_A[55]), .in_B(in_B[55]), .in_CI(1'b1), .out_S(nS_st1_b55_c1), .out_CO(nC_st1_b55_c1));
  VHA U_st1_b56_c0 (.in_A(in_A[56]), .in_B(in_B[56]), .out_S(nS_st1_b56_c0), .out_CO(nC_st1_b56_c0));
  VFA U_st1_b56_c1 (.in_A(in_A[56]), .in_B(in_B[56]), .in_CI(1'b1), .out_S(nS_st1_b56_c1), .out_CO(nC_st1_b56_c1));
  VHA U_st1_b57_c0 (.in_A(in_A[57]), .in_B(in_B[57]), .out_S(nS_st1_b57_c0), .out_CO(nC_st1_b57_c0));
  VFA U_st1_b57_c1 (.in_A(in_A[57]), .in_B(in_B[57]), .in_CI(1'b1), .out_S(nS_st1_b57_c1), .out_CO(nC_st1_b57_c1));
  VHA U_st1_b58_c0 (.in_A(in_A[58]), .in_B(in_B[58]), .out_S(nS_st1_b58_c0), .out_CO(nC_st1_b58_c0));
  VFA U_st1_b58_c1 (.in_A(in_A[58]), .in_B(in_B[58]), .in_CI(1'b1), .out_S(nS_st1_b58_c1), .out_CO(nC_st1_b58_c1));
  VHA U_st1_b59_c0 (.in_A(in_A[59]), .in_B(in_B[59]), .out_S(nS_st1_b59_c0), .out_CO(nC_st1_b59_c0));
  VFA U_st1_b59_c1 (.in_A(in_A[59]), .in_B(in_B[59]), .in_CI(1'b1), .out_S(nS_st1_b59_c1), .out_CO(nC_st1_b59_c1));
  VHA U_st1_b60_c0 (.in_A(in_A[60]), .in_B(in_B[60]), .out_S(nS_st1_b60_c0), .out_CO(nC_st1_b60_c0));
  VFA U_st1_b60_c1 (.in_A(in_A[60]), .in_B(in_B[60]), .in_CI(1'b1), .out_S(nS_st1_b60_c1), .out_CO(nC_st1_b60_c1));
  VHA U_st1_b61_c0 (.in_A(in_A[61]), .in_B(in_B[61]), .out_S(nS_st1_b61_c0), .out_CO(nC_st1_b61_c0));
  VFA U_st1_b61_c1 (.in_A(in_A[61]), .in_B(in_B[61]), .in_CI(1'b1), .out_S(nS_st1_b61_c1), .out_CO(nC_st1_b61_c1));
  VHA U_st1_b62_c0 (.in_A(in_A[62]), .in_B(in_B[62]), .out_S(nS_st1_b62_c0), .out_CO(nC_st1_b62_c0));
  VFA U_st1_b62_c1 (.in_A(in_A[62]), .in_B(in_B[62]), .in_CI(1'b1), .out_S(nS_st1_b62_c1), .out_CO(nC_st1_b62_c1));
  VHA U_st1_b63_c0 (.in_A(in_A[63]), .in_B(in_B[63]), .out_S(nS_st1_b63_c0), .out_CO(nC_st1_b63_c0));
  VFA U_st1_b63_c1 (.in_A(in_A[63]), .in_B(in_B[63]), .in_CI(1'b1), .out_S(nS_st1_b63_c1), .out_CO(nC_st1_b63_c1));
  VHA U_st1_b64_c0 (.in_A(in_A[64]), .in_B(in_B[64]), .out_S(nS_st1_b64_c0), .out_CO(nC_st1_b64_c0));
  VFA U_st1_b64_c1 (.in_A(in_A[64]), .in_B(in_B[64]), .in_CI(1'b1), .out_S(nS_st1_b64_c1), .out_CO(nC_st1_b64_c1));
  VHA U_st1_b65_c0 (.in_A(in_A[65]), .in_B(in_B[65]), .out_S(nS_st1_b65_c0), .out_CO(nC_st1_b65_c0));
  VFA U_st1_b65_c1 (.in_A(in_A[65]), .in_B(in_B[65]), .in_CI(1'b1), .out_S(nS_st1_b65_c1), .out_CO(nC_st1_b65_c1));
  VHA U_st1_b66_c0 (.in_A(in_A[66]), .in_B(in_B[66]), .out_S(nS_st1_b66_c0), .out_CO(nC_st1_b66_c0));
  VFA U_st1_b66_c1 (.in_A(in_A[66]), .in_B(in_B[66]), .in_CI(1'b1), .out_S(nS_st1_b66_c1), .out_CO(nC_st1_b66_c1));
  VHA U_st1_b67_c0 (.in_A(in_A[67]), .in_B(in_B[67]), .out_S(nS_st1_b67_c0), .out_CO(nC_st1_b67_c0));
  VFA U_st1_b67_c1 (.in_A(in_A[67]), .in_B(in_B[67]), .in_CI(1'b1), .out_S(nS_st1_b67_c1), .out_CO(nC_st1_b67_c1));
  VHA U_st1_b68_c0 (.in_A(in_A[68]), .in_B(in_B[68]), .out_S(nS_st1_b68_c0), .out_CO(nC_st1_b68_c0));
  VFA U_st1_b68_c1 (.in_A(in_A[68]), .in_B(in_B[68]), .in_CI(1'b1), .out_S(nS_st1_b68_c1), .out_CO(nC_st1_b68_c1));
  VHA U_st1_b69_c0 (.in_A(in_A[69]), .in_B(in_B[69]), .out_S(nS_st1_b69_c0), .out_CO(nC_st1_b69_c0));
  VFA U_st1_b69_c1 (.in_A(in_A[69]), .in_B(in_B[69]), .in_CI(1'b1), .out_S(nS_st1_b69_c1), .out_CO(nC_st1_b69_c1));
  VHA U_st1_b70_c0 (.in_A(in_A[70]), .in_B(in_B[70]), .out_S(nS_st1_b70_c0), .out_CO(nC_st1_b70_c0));
  VFA U_st1_b70_c1 (.in_A(in_A[70]), .in_B(in_B[70]), .in_CI(1'b1), .out_S(nS_st1_b70_c1), .out_CO(nC_st1_b70_c1));
  VHA U_st1_b71_c0 (.in_A(in_A[71]), .in_B(in_B[71]), .out_S(nS_st1_b71_c0), .out_CO(nC_st1_b71_c0));
  VFA U_st1_b71_c1 (.in_A(in_A[71]), .in_B(in_B[71]), .in_CI(1'b1), .out_S(nS_st1_b71_c1), .out_CO(nC_st1_b71_c1));
  VHA U_st1_b72_c0 (.in_A(in_A[72]), .in_B(in_B[72]), .out_S(nS_st1_b72_c0), .out_CO(nC_st1_b72_c0));
  VFA U_st1_b72_c1 (.in_A(in_A[72]), .in_B(in_B[72]), .in_CI(1'b1), .out_S(nS_st1_b72_c1), .out_CO(nC_st1_b72_c1));
  VHA U_st1_b73_c0 (.in_A(in_A[73]), .in_B(in_B[73]), .out_S(nS_st1_b73_c0), .out_CO(nC_st1_b73_c0));
  VFA U_st1_b73_c1 (.in_A(in_A[73]), .in_B(in_B[73]), .in_CI(1'b1), .out_S(nS_st1_b73_c1), .out_CO(nC_st1_b73_c1));
  VHA U_st1_b74_c0 (.in_A(in_A[74]), .in_B(in_B[74]), .out_S(nS_st1_b74_c0), .out_CO(nC_st1_b74_c0));
  VFA U_st1_b74_c1 (.in_A(in_A[74]), .in_B(in_B[74]), .in_CI(1'b1), .out_S(nS_st1_b74_c1), .out_CO(nC_st1_b74_c1));
  VHA U_st1_b75_c0 (.in_A(in_A[75]), .in_B(in_B[75]), .out_S(nS_st1_b75_c0), .out_CO(nC_st1_b75_c0));
  VFA U_st1_b75_c1 (.in_A(in_A[75]), .in_B(in_B[75]), .in_CI(1'b1), .out_S(nS_st1_b75_c1), .out_CO(nC_st1_b75_c1));
  VHA U_st1_b76_c0 (.in_A(in_A[76]), .in_B(in_B[76]), .out_S(nS_st1_b76_c0), .out_CO(nC_st1_b76_c0));
  VFA U_st1_b76_c1 (.in_A(in_A[76]), .in_B(in_B[76]), .in_CI(1'b1), .out_S(nS_st1_b76_c1), .out_CO(nC_st1_b76_c1));
  VHA U_st1_b77_c0 (.in_A(in_A[77]), .in_B(in_B[77]), .out_S(nS_st1_b77_c0), .out_CO(nC_st1_b77_c0));
  VFA U_st1_b77_c1 (.in_A(in_A[77]), .in_B(in_B[77]), .in_CI(1'b1), .out_S(nS_st1_b77_c1), .out_CO(nC_st1_b77_c1));
  VHA U_st1_b78_c0 (.in_A(in_A[78]), .in_B(in_B[78]), .out_S(nS_st1_b78_c0), .out_CO(nC_st1_b78_c0));
  VFA U_st1_b78_c1 (.in_A(in_A[78]), .in_B(in_B[78]), .in_CI(1'b1), .out_S(nS_st1_b78_c1), .out_CO(nC_st1_b78_c1));
  VHA U_st1_b79_c0 (.in_A(in_A[79]), .in_B(in_B[79]), .out_S(nS_st1_b79_c0), .out_CO(nC_st1_b79_c0));
  VFA U_st1_b79_c1 (.in_A(in_A[79]), .in_B(in_B[79]), .in_CI(1'b1), .out_S(nS_st1_b79_c1), .out_CO(nC_st1_b79_c1));
  VHA U_st1_b80_c0 (.in_A(in_A[80]), .in_B(in_B[80]), .out_S(nS_st1_b80_c0), .out_CO(nC_st1_b80_c0));
  VFA U_st1_b80_c1 (.in_A(in_A[80]), .in_B(in_B[80]), .in_CI(1'b1), .out_S(nS_st1_b80_c1), .out_CO(nC_st1_b80_c1));
  VHA U_st1_b81_c0 (.in_A(in_A[81]), .in_B(in_B[81]), .out_S(nS_st1_b81_c0), .out_CO(nC_st1_b81_c0));
  VFA U_st1_b81_c1 (.in_A(in_A[81]), .in_B(in_B[81]), .in_CI(1'b1), .out_S(nS_st1_b81_c1), .out_CO(nC_st1_b81_c1));
  VHA U_st1_b82_c0 (.in_A(in_A[82]), .in_B(in_B[82]), .out_S(nS_st1_b82_c0), .out_CO(nC_st1_b82_c0));
  VFA U_st1_b82_c1 (.in_A(in_A[82]), .in_B(in_B[82]), .in_CI(1'b1), .out_S(nS_st1_b82_c1), .out_CO(nC_st1_b82_c1));
  VHA U_st1_b83_c0 (.in_A(in_A[83]), .in_B(in_B[83]), .out_S(nS_st1_b83_c0), .out_CO(nC_st1_b83_c0));
  VFA U_st1_b83_c1 (.in_A(in_A[83]), .in_B(in_B[83]), .in_CI(1'b1), .out_S(nS_st1_b83_c1), .out_CO(nC_st1_b83_c1));
  VHA U_st1_b84_c0 (.in_A(in_A[84]), .in_B(in_B[84]), .out_S(nS_st1_b84_c0), .out_CO(nC_st1_b84_c0));
  VFA U_st1_b84_c1 (.in_A(in_A[84]), .in_B(in_B[84]), .in_CI(1'b1), .out_S(nS_st1_b84_c1), .out_CO(nC_st1_b84_c1));
  VHA U_st1_b85_c0 (.in_A(in_A[85]), .in_B(in_B[85]), .out_S(nS_st1_b85_c0), .out_CO(nC_st1_b85_c0));
  VFA U_st1_b85_c1 (.in_A(in_A[85]), .in_B(in_B[85]), .in_CI(1'b1), .out_S(nS_st1_b85_c1), .out_CO(nC_st1_b85_c1));
  VHA U_st1_b86_c0 (.in_A(in_A[86]), .in_B(in_B[86]), .out_S(nS_st1_b86_c0), .out_CO(nC_st1_b86_c0));
  VFA U_st1_b86_c1 (.in_A(in_A[86]), .in_B(in_B[86]), .in_CI(1'b1), .out_S(nS_st1_b86_c1), .out_CO(nC_st1_b86_c1));
  VHA U_st1_b87_c0 (.in_A(in_A[87]), .in_B(in_B[87]), .out_S(nS_st1_b87_c0), .out_CO(nC_st1_b87_c0));
  VFA U_st1_b87_c1 (.in_A(in_A[87]), .in_B(in_B[87]), .in_CI(1'b1), .out_S(nS_st1_b87_c1), .out_CO(nC_st1_b87_c1));
  VHA U_st1_b88_c0 (.in_A(in_A[88]), .in_B(in_B[88]), .out_S(nS_st1_b88_c0), .out_CO(nC_st1_b88_c0));
  VFA U_st1_b88_c1 (.in_A(in_A[88]), .in_B(in_B[88]), .in_CI(1'b1), .out_S(nS_st1_b88_c1), .out_CO(nC_st1_b88_c1));
  VHA U_st1_b89_c0 (.in_A(in_A[89]), .in_B(in_B[89]), .out_S(nS_st1_b89_c0), .out_CO(nC_st1_b89_c0));
  VFA U_st1_b89_c1 (.in_A(in_A[89]), .in_B(in_B[89]), .in_CI(1'b1), .out_S(nS_st1_b89_c1), .out_CO(nC_st1_b89_c1));
  VHA U_st1_b90_c0 (.in_A(in_A[90]), .in_B(in_B[90]), .out_S(nS_st1_b90_c0), .out_CO(nC_st1_b90_c0));
  VFA U_st1_b90_c1 (.in_A(in_A[90]), .in_B(in_B[90]), .in_CI(1'b1), .out_S(nS_st1_b90_c1), .out_CO(nC_st1_b90_c1));
  VHA U_st1_b91_c0 (.in_A(in_A[91]), .in_B(in_B[91]), .out_S(nS_st1_b91_c0), .out_CO(nC_st1_b91_c0));
  VFA U_st1_b91_c1 (.in_A(in_A[91]), .in_B(in_B[91]), .in_CI(1'b1), .out_S(nS_st1_b91_c1), .out_CO(nC_st1_b91_c1));
  VHA U_st1_b92_c0 (.in_A(in_A[92]), .in_B(in_B[92]), .out_S(nS_st1_b92_c0), .out_CO(nC_st1_b92_c0));
  VFA U_st1_b92_c1 (.in_A(in_A[92]), .in_B(in_B[92]), .in_CI(1'b1), .out_S(nS_st1_b92_c1), .out_CO(nC_st1_b92_c1));
  VHA U_st1_b93_c0 (.in_A(in_A[93]), .in_B(in_B[93]), .out_S(nS_st1_b93_c0), .out_CO(nC_st1_b93_c0));
  VFA U_st1_b93_c1 (.in_A(in_A[93]), .in_B(in_B[93]), .in_CI(1'b1), .out_S(nS_st1_b93_c1), .out_CO(nC_st1_b93_c1));
  VHA U_st1_b94_c0 (.in_A(in_A[94]), .in_B(in_B[94]), .out_S(nS_st1_b94_c0), .out_CO(nC_st1_b94_c0));
  VFA U_st1_b94_c1 (.in_A(in_A[94]), .in_B(in_B[94]), .in_CI(1'b1), .out_S(nS_st1_b94_c1), .out_CO(nC_st1_b94_c1));
  VHA U_st1_b95_c0 (.in_A(in_A[95]), .in_B(in_B[95]), .out_S(nS_st1_b95_c0), .out_CO(nC_st1_b95_c0));
  VFA U_st1_b95_c1 (.in_A(in_A[95]), .in_B(in_B[95]), .in_CI(1'b1), .out_S(nS_st1_b95_c1), .out_CO(nC_st1_b95_c1));
  VHA U_st1_b96_c0 (.in_A(in_A[96]), .in_B(in_B[96]), .out_S(nS_st1_b96_c0), .out_CO(nC_st1_b96_c0));
  VFA U_st1_b96_c1 (.in_A(in_A[96]), .in_B(in_B[96]), .in_CI(1'b1), .out_S(nS_st1_b96_c1), .out_CO(nC_st1_b96_c1));
  VHA U_st1_b97_c0 (.in_A(in_A[97]), .in_B(in_B[97]), .out_S(nS_st1_b97_c0), .out_CO(nC_st1_b97_c0));
  VFA U_st1_b97_c1 (.in_A(in_A[97]), .in_B(in_B[97]), .in_CI(1'b1), .out_S(nS_st1_b97_c1), .out_CO(nC_st1_b97_c1));
  VHA U_st1_b98_c0 (.in_A(in_A[98]), .in_B(in_B[98]), .out_S(nS_st1_b98_c0), .out_CO(nC_st1_b98_c0));
  VFA U_st1_b98_c1 (.in_A(in_A[98]), .in_B(in_B[98]), .in_CI(1'b1), .out_S(nS_st1_b98_c1), .out_CO(nC_st1_b98_c1));
  VHA U_st1_b99_c0 (.in_A(in_A[99]), .in_B(in_B[99]), .out_S(nS_st1_b99_c0), .out_CO(nC_st1_b99_c0));
  VFA U_st1_b99_c1 (.in_A(in_A[99]), .in_B(in_B[99]), .in_CI(1'b1), .out_S(nS_st1_b99_c1), .out_CO(nC_st1_b99_c1));
  VHA U_st1_b100_c0 (.in_A(in_A[100]), .in_B(in_B[100]), .out_S(nS_st1_b100_c0), .out_CO(nC_st1_b100_c0));
  VFA U_st1_b100_c1 (.in_A(in_A[100]), .in_B(in_B[100]), .in_CI(1'b1), .out_S(nS_st1_b100_c1), .out_CO(nC_st1_b100_c1));
  VHA U_st1_b101_c0 (.in_A(in_A[101]), .in_B(in_B[101]), .out_S(nS_st1_b101_c0), .out_CO(nC_st1_b101_c0));
  VFA U_st1_b101_c1 (.in_A(in_A[101]), .in_B(in_B[101]), .in_CI(1'b1), .out_S(nS_st1_b101_c1), .out_CO(nC_st1_b101_c1));
  VHA U_st1_b102_c0 (.in_A(in_A[102]), .in_B(in_B[102]), .out_S(nS_st1_b102_c0), .out_CO(nC_st1_b102_c0));
  VFA U_st1_b102_c1 (.in_A(in_A[102]), .in_B(in_B[102]), .in_CI(1'b1), .out_S(nS_st1_b102_c1), .out_CO(nC_st1_b102_c1));
  VHA U_st1_b103_c0 (.in_A(in_A[103]), .in_B(in_B[103]), .out_S(nS_st1_b103_c0), .out_CO(nC_st1_b103_c0));
  VFA U_st1_b103_c1 (.in_A(in_A[103]), .in_B(in_B[103]), .in_CI(1'b1), .out_S(nS_st1_b103_c1), .out_CO(nC_st1_b103_c1));
  VHA U_st1_b104_c0 (.in_A(in_A[104]), .in_B(in_B[104]), .out_S(nS_st1_b104_c0), .out_CO(nC_st1_b104_c0));
  VFA U_st1_b104_c1 (.in_A(in_A[104]), .in_B(in_B[104]), .in_CI(1'b1), .out_S(nS_st1_b104_c1), .out_CO(nC_st1_b104_c1));
  VHA U_st1_b105_c0 (.in_A(in_A[105]), .in_B(in_B[105]), .out_S(nS_st1_b105_c0), .out_CO(nC_st1_b105_c0));
  VFA U_st1_b105_c1 (.in_A(in_A[105]), .in_B(in_B[105]), .in_CI(1'b1), .out_S(nS_st1_b105_c1), .out_CO(nC_st1_b105_c1));
  VHA U_st1_b106_c0 (.in_A(in_A[106]), .in_B(in_B[106]), .out_S(nS_st1_b106_c0), .out_CO(nC_st1_b106_c0));
  VFA U_st1_b106_c1 (.in_A(in_A[106]), .in_B(in_B[106]), .in_CI(1'b1), .out_S(nS_st1_b106_c1), .out_CO(nC_st1_b106_c1));
  VHA U_st1_b107_c0 (.in_A(in_A[107]), .in_B(in_B[107]), .out_S(nS_st1_b107_c0), .out_CO(nC_st1_b107_c0));
  VFA U_st1_b107_c1 (.in_A(in_A[107]), .in_B(in_B[107]), .in_CI(1'b1), .out_S(nS_st1_b107_c1), .out_CO(nC_st1_b107_c1));
  VHA U_st1_b108_c0 (.in_A(in_A[108]), .in_B(in_B[108]), .out_S(nS_st1_b108_c0), .out_CO(nC_st1_b108_c0));
  VFA U_st1_b108_c1 (.in_A(in_A[108]), .in_B(in_B[108]), .in_CI(1'b1), .out_S(nS_st1_b108_c1), .out_CO(nC_st1_b108_c1));
  VHA U_st1_b109_c0 (.in_A(in_A[109]), .in_B(in_B[109]), .out_S(nS_st1_b109_c0), .out_CO(nC_st1_b109_c0));
  VFA U_st1_b109_c1 (.in_A(in_A[109]), .in_B(in_B[109]), .in_CI(1'b1), .out_S(nS_st1_b109_c1), .out_CO(nC_st1_b109_c1));
  VHA U_st1_b110_c0 (.in_A(in_A[110]), .in_B(in_B[110]), .out_S(nS_st1_b110_c0), .out_CO(nC_st1_b110_c0));
  VFA U_st1_b110_c1 (.in_A(in_A[110]), .in_B(in_B[110]), .in_CI(1'b1), .out_S(nS_st1_b110_c1), .out_CO(nC_st1_b110_c1));
  VHA U_st1_b111_c0 (.in_A(in_A[111]), .in_B(in_B[111]), .out_S(nS_st1_b111_c0), .out_CO(nC_st1_b111_c0));
  VFA U_st1_b111_c1 (.in_A(in_A[111]), .in_B(in_B[111]), .in_CI(1'b1), .out_S(nS_st1_b111_c1), .out_CO(nC_st1_b111_c1));
  VHA U_st1_b112_c0 (.in_A(in_A[112]), .in_B(in_B[112]), .out_S(nS_st1_b112_c0), .out_CO(nC_st1_b112_c0));
  VFA U_st1_b112_c1 (.in_A(in_A[112]), .in_B(in_B[112]), .in_CI(1'b1), .out_S(nS_st1_b112_c1), .out_CO(nC_st1_b112_c1));
  VHA U_st1_b113_c0 (.in_A(in_A[113]), .in_B(in_B[113]), .out_S(nS_st1_b113_c0), .out_CO(nC_st1_b113_c0));
  VFA U_st1_b113_c1 (.in_A(in_A[113]), .in_B(in_B[113]), .in_CI(1'b1), .out_S(nS_st1_b113_c1), .out_CO(nC_st1_b113_c1));
  VHA U_st1_b114_c0 (.in_A(in_A[114]), .in_B(in_B[114]), .out_S(nS_st1_b114_c0), .out_CO(nC_st1_b114_c0));
  VFA U_st1_b114_c1 (.in_A(in_A[114]), .in_B(in_B[114]), .in_CI(1'b1), .out_S(nS_st1_b114_c1), .out_CO(nC_st1_b114_c1));
  VHA U_st1_b115_c0 (.in_A(in_A[115]), .in_B(in_B[115]), .out_S(nS_st1_b115_c0), .out_CO(nC_st1_b115_c0));
  VFA U_st1_b115_c1 (.in_A(in_A[115]), .in_B(in_B[115]), .in_CI(1'b1), .out_S(nS_st1_b115_c1), .out_CO(nC_st1_b115_c1));
  VHA U_st1_b116_c0 (.in_A(in_A[116]), .in_B(in_B[116]), .out_S(nS_st1_b116_c0), .out_CO(nC_st1_b116_c0));
  VFA U_st1_b116_c1 (.in_A(in_A[116]), .in_B(in_B[116]), .in_CI(1'b1), .out_S(nS_st1_b116_c1), .out_CO(nC_st1_b116_c1));
  VHA U_st1_b117_c0 (.in_A(in_A[117]), .in_B(in_B[117]), .out_S(nS_st1_b117_c0), .out_CO(nC_st1_b117_c0));
  VFA U_st1_b117_c1 (.in_A(in_A[117]), .in_B(in_B[117]), .in_CI(1'b1), .out_S(nS_st1_b117_c1), .out_CO(nC_st1_b117_c1));
  VHA U_st1_b118_c0 (.in_A(in_A[118]), .in_B(in_B[118]), .out_S(nS_st1_b118_c0), .out_CO(nC_st1_b118_c0));
  VFA U_st1_b118_c1 (.in_A(in_A[118]), .in_B(in_B[118]), .in_CI(1'b1), .out_S(nS_st1_b118_c1), .out_CO(nC_st1_b118_c1));
  VHA U_st1_b119_c0 (.in_A(in_A[119]), .in_B(in_B[119]), .out_S(nS_st1_b119_c0), .out_CO(nC_st1_b119_c0));
  VFA U_st1_b119_c1 (.in_A(in_A[119]), .in_B(in_B[119]), .in_CI(1'b1), .out_S(nS_st1_b119_c1), .out_CO(nC_st1_b119_c1));
  VHA U_st1_b120_c0 (.in_A(in_A[120]), .in_B(in_B[120]), .out_S(nS_st1_b120_c0), .out_CO(nC_st1_b120_c0));
  VFA U_st1_b120_c1 (.in_A(in_A[120]), .in_B(in_B[120]), .in_CI(1'b1), .out_S(nS_st1_b120_c1), .out_CO(nC_st1_b120_c1));
  VHA U_st1_b121_c0 (.in_A(in_A[121]), .in_B(in_B[121]), .out_S(nS_st1_b121_c0), .out_CO(nC_st1_b121_c0));
  VFA U_st1_b121_c1 (.in_A(in_A[121]), .in_B(in_B[121]), .in_CI(1'b1), .out_S(nS_st1_b121_c1), .out_CO(nC_st1_b121_c1));
  VHA U_st1_b122_c0 (.in_A(in_A[122]), .in_B(in_B[122]), .out_S(nS_st1_b122_c0), .out_CO(nC_st1_b122_c0));
  VFA U_st1_b122_c1 (.in_A(in_A[122]), .in_B(in_B[122]), .in_CI(1'b1), .out_S(nS_st1_b122_c1), .out_CO(nC_st1_b122_c1));
  VHA U_st1_b123_c0 (.in_A(in_A[123]), .in_B(in_B[123]), .out_S(nS_st1_b123_c0), .out_CO(nC_st1_b123_c0));
  VFA U_st1_b123_c1 (.in_A(in_A[123]), .in_B(in_B[123]), .in_CI(1'b1), .out_S(nS_st1_b123_c1), .out_CO(nC_st1_b123_c1));
  VHA U_st1_b124_c0 (.in_A(in_A[124]), .in_B(in_B[124]), .out_S(nS_st1_b124_c0), .out_CO(nC_st1_b124_c0));
  VFA U_st1_b124_c1 (.in_A(in_A[124]), .in_B(in_B[124]), .in_CI(1'b1), .out_S(nS_st1_b124_c1), .out_CO(nC_st1_b124_c1));
  VHA U_st1_b125_c0 (.in_A(in_A[125]), .in_B(in_B[125]), .out_S(nS_st1_b125_c0), .out_CO(nC_st1_b125_c0));
  VFA U_st1_b125_c1 (.in_A(in_A[125]), .in_B(in_B[125]), .in_CI(1'b1), .out_S(nS_st1_b125_c1), .out_CO(nC_st1_b125_c1));
  VHA U_st1_b126_c0 (.in_A(in_A[126]), .in_B(in_B[126]), .out_S(nS_st1_b126_c0), .out_CO(nC_st1_b126_c0));
  VFA U_st1_b126_c1 (.in_A(in_A[126]), .in_B(in_B[126]), .in_CI(1'b1), .out_S(nS_st1_b126_c1), .out_CO(nC_st1_b126_c1));
  VHA U_st1_b127_c0 (.in_A(in_A[127]), .in_B(in_B[127]), .out_S(nS_st1_b127_c0), .out_CO(nC_st1_b127_c0));
  VFA U_st1_b127_c1 (.in_A(in_A[127]), .in_B(in_B[127]), .in_CI(1'b1), .out_S(nS_st1_b127_c1), .out_CO(nC_st1_b127_c1));
  VHA U_st1_b128_c0 (.in_A(in_A[128]), .in_B(in_B[128]), .out_S(nS_st1_b128_c0), .out_CO(nC_st1_b128_c0));
  VFA U_st1_b128_c1 (.in_A(in_A[128]), .in_B(in_B[128]), .in_CI(1'b1), .out_S(nS_st1_b128_c1), .out_CO(nC_st1_b128_c1));
  VHA U_st1_b129_c0 (.in_A(in_A[129]), .in_B(in_B[129]), .out_S(nS_st1_b129_c0), .out_CO(nC_st1_b129_c0));
  VFA U_st1_b129_c1 (.in_A(in_A[129]), .in_B(in_B[129]), .in_CI(1'b1), .out_S(nS_st1_b129_c1), .out_CO(nC_st1_b129_c1));
  VHA U_st1_b130_c0 (.in_A(in_A[130]), .in_B(in_B[130]), .out_S(nS_st1_b130_c0), .out_CO(nC_st1_b130_c0));
  VFA U_st1_b130_c1 (.in_A(in_A[130]), .in_B(in_B[130]), .in_CI(1'b1), .out_S(nS_st1_b130_c1), .out_CO(nC_st1_b130_c1));
  VHA U_st1_b131_c0 (.in_A(in_A[131]), .in_B(in_B[131]), .out_S(nS_st1_b131_c0), .out_CO(nC_st1_b131_c0));
  VFA U_st1_b131_c1 (.in_A(in_A[131]), .in_B(in_B[131]), .in_CI(1'b1), .out_S(nS_st1_b131_c1), .out_CO(nC_st1_b131_c1));
  VHA U_st1_b132_c0 (.in_A(in_A[132]), .in_B(in_B[132]), .out_S(nS_st1_b132_c0), .out_CO(nC_st1_b132_c0));
  VFA U_st1_b132_c1 (.in_A(in_A[132]), .in_B(in_B[132]), .in_CI(1'b1), .out_S(nS_st1_b132_c1), .out_CO(nC_st1_b132_c1));
  VHA U_st1_b133_c0 (.in_A(in_A[133]), .in_B(in_B[133]), .out_S(nS_st1_b133_c0), .out_CO(nC_st1_b133_c0));
  VFA U_st1_b133_c1 (.in_A(in_A[133]), .in_B(in_B[133]), .in_CI(1'b1), .out_S(nS_st1_b133_c1), .out_CO(nC_st1_b133_c1));
  VHA U_st1_b134_c0 (.in_A(in_A[134]), .in_B(in_B[134]), .out_S(nS_st1_b134_c0), .out_CO(nC_st1_b134_c0));
  VFA U_st1_b134_c1 (.in_A(in_A[134]), .in_B(in_B[134]), .in_CI(1'b1), .out_S(nS_st1_b134_c1), .out_CO(nC_st1_b134_c1));
  VHA U_st1_b135_c0 (.in_A(in_A[135]), .in_B(in_B[135]), .out_S(nS_st1_b135_c0), .out_CO(nC_st1_b135_c0));
  VFA U_st1_b135_c1 (.in_A(in_A[135]), .in_B(in_B[135]), .in_CI(1'b1), .out_S(nS_st1_b135_c1), .out_CO(nC_st1_b135_c1));
  VHA U_st1_b136_c0 (.in_A(in_A[136]), .in_B(in_B[136]), .out_S(nS_st1_b136_c0), .out_CO(nC_st1_b136_c0));
  VFA U_st1_b136_c1 (.in_A(in_A[136]), .in_B(in_B[136]), .in_CI(1'b1), .out_S(nS_st1_b136_c1), .out_CO(nC_st1_b136_c1));
  VHA U_st1_b137_c0 (.in_A(in_A[137]), .in_B(in_B[137]), .out_S(nS_st1_b137_c0), .out_CO(nC_st1_b137_c0));
  VFA U_st1_b137_c1 (.in_A(in_A[137]), .in_B(in_B[137]), .in_CI(1'b1), .out_S(nS_st1_b137_c1), .out_CO(nC_st1_b137_c1));
  VHA U_st1_b138_c0 (.in_A(in_A[138]), .in_B(in_B[138]), .out_S(nS_st1_b138_c0), .out_CO(nC_st1_b138_c0));
  VFA U_st1_b138_c1 (.in_A(in_A[138]), .in_B(in_B[138]), .in_CI(1'b1), .out_S(nS_st1_b138_c1), .out_CO(nC_st1_b138_c1));
  VHA U_st1_b139_c0 (.in_A(in_A[139]), .in_B(in_B[139]), .out_S(nS_st1_b139_c0), .out_CO(nC_st1_b139_c0));
  VFA U_st1_b139_c1 (.in_A(in_A[139]), .in_B(in_B[139]), .in_CI(1'b1), .out_S(nS_st1_b139_c1), .out_CO(nC_st1_b139_c1));
  VHA U_st1_b140_c0 (.in_A(in_A[140]), .in_B(in_B[140]), .out_S(nS_st1_b140_c0), .out_CO(nC_st1_b140_c0));
  VFA U_st1_b140_c1 (.in_A(in_A[140]), .in_B(in_B[140]), .in_CI(1'b1), .out_S(nS_st1_b140_c1), .out_CO(nC_st1_b140_c1));
  VHA U_st1_b141_c0 (.in_A(in_A[141]), .in_B(in_B[141]), .out_S(nS_st1_b141_c0), .out_CO(nC_st1_b141_c0));
  VFA U_st1_b141_c1 (.in_A(in_A[141]), .in_B(in_B[141]), .in_CI(1'b1), .out_S(nS_st1_b141_c1), .out_CO(nC_st1_b141_c1));
  VHA U_st1_b142_c0 (.in_A(in_A[142]), .in_B(in_B[142]), .out_S(nS_st1_b142_c0), .out_CO(nC_st1_b142_c0));
  VFA U_st1_b142_c1 (.in_A(in_A[142]), .in_B(in_B[142]), .in_CI(1'b1), .out_S(nS_st1_b142_c1), .out_CO(nC_st1_b142_c1));
  VHA U_st1_b143_c0 (.in_A(in_A[143]), .in_B(in_B[143]), .out_S(nS_st1_b143_c0), .out_CO(nC_st1_b143_c0));
  VFA U_st1_b143_c1 (.in_A(in_A[143]), .in_B(in_B[143]), .in_CI(1'b1), .out_S(nS_st1_b143_c1), .out_CO(nC_st1_b143_c1));
  VHA U_st1_b144_c0 (.in_A(in_A[144]), .in_B(in_B[144]), .out_S(nS_st1_b144_c0), .out_CO(nC_st1_b144_c0));
  VFA U_st1_b144_c1 (.in_A(in_A[144]), .in_B(in_B[144]), .in_CI(1'b1), .out_S(nS_st1_b144_c1), .out_CO(nC_st1_b144_c1));
  VHA U_st1_b145_c0 (.in_A(in_A[145]), .in_B(in_B[145]), .out_S(nS_st1_b145_c0), .out_CO(nC_st1_b145_c0));
  VFA U_st1_b145_c1 (.in_A(in_A[145]), .in_B(in_B[145]), .in_CI(1'b1), .out_S(nS_st1_b145_c1), .out_CO(nC_st1_b145_c1));
  VHA U_st1_b146_c0 (.in_A(in_A[146]), .in_B(in_B[146]), .out_S(nS_st1_b146_c0), .out_CO(nC_st1_b146_c0));
  VFA U_st1_b146_c1 (.in_A(in_A[146]), .in_B(in_B[146]), .in_CI(1'b1), .out_S(nS_st1_b146_c1), .out_CO(nC_st1_b146_c1));
  VHA U_st1_b147_c0 (.in_A(in_A[147]), .in_B(in_B[147]), .out_S(nS_st1_b147_c0), .out_CO(nC_st1_b147_c0));
  VFA U_st1_b147_c1 (.in_A(in_A[147]), .in_B(in_B[147]), .in_CI(1'b1), .out_S(nS_st1_b147_c1), .out_CO(nC_st1_b147_c1));
  VHA U_st1_b148_c0 (.in_A(in_A[148]), .in_B(in_B[148]), .out_S(nS_st1_b148_c0), .out_CO(nC_st1_b148_c0));
  VFA U_st1_b148_c1 (.in_A(in_A[148]), .in_B(in_B[148]), .in_CI(1'b1), .out_S(nS_st1_b148_c1), .out_CO(nC_st1_b148_c1));
  VHA U_st1_b149_c0 (.in_A(in_A[149]), .in_B(in_B[149]), .out_S(nS_st1_b149_c0), .out_CO(nC_st1_b149_c0));
  VFA U_st1_b149_c1 (.in_A(in_A[149]), .in_B(in_B[149]), .in_CI(1'b1), .out_S(nS_st1_b149_c1), .out_CO(nC_st1_b149_c1));
  VHA U_st1_b150_c0 (.in_A(in_A[150]), .in_B(in_B[150]), .out_S(nS_st1_b150_c0), .out_CO(nC_st1_b150_c0));
  VFA U_st1_b150_c1 (.in_A(in_A[150]), .in_B(in_B[150]), .in_CI(1'b1), .out_S(nS_st1_b150_c1), .out_CO(nC_st1_b150_c1));
  VHA U_st1_b151_c0 (.in_A(in_A[151]), .in_B(in_B[151]), .out_S(nS_st1_b151_c0), .out_CO(nC_st1_b151_c0));
  VFA U_st1_b151_c1 (.in_A(in_A[151]), .in_B(in_B[151]), .in_CI(1'b1), .out_S(nS_st1_b151_c1), .out_CO(nC_st1_b151_c1));
  VHA U_st1_b152_c0 (.in_A(in_A[152]), .in_B(in_B[152]), .out_S(nS_st1_b152_c0), .out_CO(nC_st1_b152_c0));
  VFA U_st1_b152_c1 (.in_A(in_A[152]), .in_B(in_B[152]), .in_CI(1'b1), .out_S(nS_st1_b152_c1), .out_CO(nC_st1_b152_c1));
  VHA U_st1_b153_c0 (.in_A(in_A[153]), .in_B(in_B[153]), .out_S(nS_st1_b153_c0), .out_CO(nC_st1_b153_c0));
  VFA U_st1_b153_c1 (.in_A(in_A[153]), .in_B(in_B[153]), .in_CI(1'b1), .out_S(nS_st1_b153_c1), .out_CO(nC_st1_b153_c1));
  VHA U_st1_b154_c0 (.in_A(in_A[154]), .in_B(in_B[154]), .out_S(nS_st1_b154_c0), .out_CO(nC_st1_b154_c0));
  VFA U_st1_b154_c1 (.in_A(in_A[154]), .in_B(in_B[154]), .in_CI(1'b1), .out_S(nS_st1_b154_c1), .out_CO(nC_st1_b154_c1));
  VHA U_st1_b155_c0 (.in_A(in_A[155]), .in_B(in_B[155]), .out_S(nS_st1_b155_c0), .out_CO(nC_st1_b155_c0));
  VFA U_st1_b155_c1 (.in_A(in_A[155]), .in_B(in_B[155]), .in_CI(1'b1), .out_S(nS_st1_b155_c1), .out_CO(nC_st1_b155_c1));
  VHA U_st1_b156_c0 (.in_A(in_A[156]), .in_B(in_B[156]), .out_S(nS_st1_b156_c0), .out_CO(nC_st1_b156_c0));
  VFA U_st1_b156_c1 (.in_A(in_A[156]), .in_B(in_B[156]), .in_CI(1'b1), .out_S(nS_st1_b156_c1), .out_CO(nC_st1_b156_c1));
  VHA U_st1_b157_c0 (.in_A(in_A[157]), .in_B(in_B[157]), .out_S(nS_st1_b157_c0), .out_CO(nC_st1_b157_c0));
  VFA U_st1_b157_c1 (.in_A(in_A[157]), .in_B(in_B[157]), .in_CI(1'b1), .out_S(nS_st1_b157_c1), .out_CO(nC_st1_b157_c1));
  VHA U_st1_b158_c0 (.in_A(in_A[158]), .in_B(in_B[158]), .out_S(nS_st1_b158_c0), .out_CO(nC_st1_b158_c0));
  VFA U_st1_b158_c1 (.in_A(in_A[158]), .in_B(in_B[158]), .in_CI(1'b1), .out_S(nS_st1_b158_c1), .out_CO(nC_st1_b158_c1));
  VHA U_st1_b159_c0 (.in_A(in_A[159]), .in_B(in_B[159]), .out_S(nS_st1_b159_c0), .out_CO(nC_st1_b159_c0));
  VFA U_st1_b159_c1 (.in_A(in_A[159]), .in_B(in_B[159]), .in_CI(1'b1), .out_S(nS_st1_b159_c1), .out_CO(nC_st1_b159_c1));
  VHA U_st1_b160_c0 (.in_A(in_A[160]), .in_B(in_B[160]), .out_S(nS_st1_b160_c0), .out_CO(nC_st1_b160_c0));
  VFA U_st1_b160_c1 (.in_A(in_A[160]), .in_B(in_B[160]), .in_CI(1'b1), .out_S(nS_st1_b160_c1), .out_CO(nC_st1_b160_c1));
  VHA U_st1_b161_c0 (.in_A(in_A[161]), .in_B(in_B[161]), .out_S(nS_st1_b161_c0), .out_CO(nC_st1_b161_c0));
  VFA U_st1_b161_c1 (.in_A(in_A[161]), .in_B(in_B[161]), .in_CI(1'b1), .out_S(nS_st1_b161_c1), .out_CO(nC_st1_b161_c1));
  VHA U_st1_b162_c0 (.in_A(in_A[162]), .in_B(in_B[162]), .out_S(nS_st1_b162_c0), .out_CO(nC_st1_b162_c0));
  VFA U_st1_b162_c1 (.in_A(in_A[162]), .in_B(in_B[162]), .in_CI(1'b1), .out_S(nS_st1_b162_c1), .out_CO(nC_st1_b162_c1));
  VHA U_st1_b163_c0 (.in_A(in_A[163]), .in_B(in_B[163]), .out_S(nS_st1_b163_c0), .out_CO(nC_st1_b163_c0));
  VFA U_st1_b163_c1 (.in_A(in_A[163]), .in_B(in_B[163]), .in_CI(1'b1), .out_S(nS_st1_b163_c1), .out_CO(nC_st1_b163_c1));
  VHA U_st1_b164_c0 (.in_A(in_A[164]), .in_B(in_B[164]), .out_S(nS_st1_b164_c0), .out_CO(nC_st1_b164_c0));
  VFA U_st1_b164_c1 (.in_A(in_A[164]), .in_B(in_B[164]), .in_CI(1'b1), .out_S(nS_st1_b164_c1), .out_CO(nC_st1_b164_c1));
  VHA U_st1_b165_c0 (.in_A(in_A[165]), .in_B(in_B[165]), .out_S(nS_st1_b165_c0), .out_CO(nC_st1_b165_c0));
  VFA U_st1_b165_c1 (.in_A(in_A[165]), .in_B(in_B[165]), .in_CI(1'b1), .out_S(nS_st1_b165_c1), .out_CO(nC_st1_b165_c1));
  VHA U_st1_b166_c0 (.in_A(in_A[166]), .in_B(in_B[166]), .out_S(nS_st1_b166_c0), .out_CO(nC_st1_b166_c0));
  VFA U_st1_b166_c1 (.in_A(in_A[166]), .in_B(in_B[166]), .in_CI(1'b1), .out_S(nS_st1_b166_c1), .out_CO(nC_st1_b166_c1));
  VHA U_st1_b167_c0 (.in_A(in_A[167]), .in_B(in_B[167]), .out_S(nS_st1_b167_c0), .out_CO(nC_st1_b167_c0));
  VFA U_st1_b167_c1 (.in_A(in_A[167]), .in_B(in_B[167]), .in_CI(1'b1), .out_S(nS_st1_b167_c1), .out_CO(nC_st1_b167_c1));
  VHA U_st1_b168_c0 (.in_A(in_A[168]), .in_B(in_B[168]), .out_S(nS_st1_b168_c0), .out_CO(nC_st1_b168_c0));
  VFA U_st1_b168_c1 (.in_A(in_A[168]), .in_B(in_B[168]), .in_CI(1'b1), .out_S(nS_st1_b168_c1), .out_CO(nC_st1_b168_c1));
  VHA U_st1_b169_c0 (.in_A(in_A[169]), .in_B(in_B[169]), .out_S(nS_st1_b169_c0), .out_CO(nC_st1_b169_c0));
  VFA U_st1_b169_c1 (.in_A(in_A[169]), .in_B(in_B[169]), .in_CI(1'b1), .out_S(nS_st1_b169_c1), .out_CO(nC_st1_b169_c1));
  VHA U_st1_b170_c0 (.in_A(in_A[170]), .in_B(in_B[170]), .out_S(nS_st1_b170_c0), .out_CO(nC_st1_b170_c0));
  VFA U_st1_b170_c1 (.in_A(in_A[170]), .in_B(in_B[170]), .in_CI(1'b1), .out_S(nS_st1_b170_c1), .out_CO(nC_st1_b170_c1));
  VHA U_st1_b171_c0 (.in_A(in_A[171]), .in_B(in_B[171]), .out_S(nS_st1_b171_c0), .out_CO(nC_st1_b171_c0));
  VFA U_st1_b171_c1 (.in_A(in_A[171]), .in_B(in_B[171]), .in_CI(1'b1), .out_S(nS_st1_b171_c1), .out_CO(nC_st1_b171_c1));
  VHA U_st1_b172_c0 (.in_A(in_A[172]), .in_B(in_B[172]), .out_S(nS_st1_b172_c0), .out_CO(nC_st1_b172_c0));
  VFA U_st1_b172_c1 (.in_A(in_A[172]), .in_B(in_B[172]), .in_CI(1'b1), .out_S(nS_st1_b172_c1), .out_CO(nC_st1_b172_c1));
  VHA U_st1_b173_c0 (.in_A(in_A[173]), .in_B(in_B[173]), .out_S(nS_st1_b173_c0), .out_CO(nC_st1_b173_c0));
  VFA U_st1_b173_c1 (.in_A(in_A[173]), .in_B(in_B[173]), .in_CI(1'b1), .out_S(nS_st1_b173_c1), .out_CO(nC_st1_b173_c1));
  VHA U_st1_b174_c0 (.in_A(in_A[174]), .in_B(in_B[174]), .out_S(nS_st1_b174_c0), .out_CO(nC_st1_b174_c0));
  VFA U_st1_b174_c1 (.in_A(in_A[174]), .in_B(in_B[174]), .in_CI(1'b1), .out_S(nS_st1_b174_c1), .out_CO(nC_st1_b174_c1));
  VHA U_st1_b175_c0 (.in_A(in_A[175]), .in_B(in_B[175]), .out_S(nS_st1_b175_c0), .out_CO(nC_st1_b175_c0));
  VFA U_st1_b175_c1 (.in_A(in_A[175]), .in_B(in_B[175]), .in_CI(1'b1), .out_S(nS_st1_b175_c1), .out_CO(nC_st1_b175_c1));
  VHA U_st1_b176_c0 (.in_A(in_A[176]), .in_B(in_B[176]), .out_S(nS_st1_b176_c0), .out_CO(nC_st1_b176_c0));
  VFA U_st1_b176_c1 (.in_A(in_A[176]), .in_B(in_B[176]), .in_CI(1'b1), .out_S(nS_st1_b176_c1), .out_CO(nC_st1_b176_c1));
  VHA U_st1_b177_c0 (.in_A(in_A[177]), .in_B(in_B[177]), .out_S(nS_st1_b177_c0), .out_CO(nC_st1_b177_c0));
  VFA U_st1_b177_c1 (.in_A(in_A[177]), .in_B(in_B[177]), .in_CI(1'b1), .out_S(nS_st1_b177_c1), .out_CO(nC_st1_b177_c1));
  VHA U_st1_b178_c0 (.in_A(in_A[178]), .in_B(in_B[178]), .out_S(nS_st1_b178_c0), .out_CO(nC_st1_b178_c0));
  VFA U_st1_b178_c1 (.in_A(in_A[178]), .in_B(in_B[178]), .in_CI(1'b1), .out_S(nS_st1_b178_c1), .out_CO(nC_st1_b178_c1));
  VHA U_st1_b179_c0 (.in_A(in_A[179]), .in_B(in_B[179]), .out_S(nS_st1_b179_c0), .out_CO(nC_st1_b179_c0));
  VFA U_st1_b179_c1 (.in_A(in_A[179]), .in_B(in_B[179]), .in_CI(1'b1), .out_S(nS_st1_b179_c1), .out_CO(nC_st1_b179_c1));
  VHA U_st1_b180_c0 (.in_A(in_A[180]), .in_B(in_B[180]), .out_S(nS_st1_b180_c0), .out_CO(nC_st1_b180_c0));
  VFA U_st1_b180_c1 (.in_A(in_A[180]), .in_B(in_B[180]), .in_CI(1'b1), .out_S(nS_st1_b180_c1), .out_CO(nC_st1_b180_c1));
  VHA U_st1_b181_c0 (.in_A(in_A[181]), .in_B(in_B[181]), .out_S(nS_st1_b181_c0), .out_CO(nC_st1_b181_c0));
  VFA U_st1_b181_c1 (.in_A(in_A[181]), .in_B(in_B[181]), .in_CI(1'b1), .out_S(nS_st1_b181_c1), .out_CO(nC_st1_b181_c1));
  VHA U_st1_b182_c0 (.in_A(in_A[182]), .in_B(in_B[182]), .out_S(nS_st1_b182_c0), .out_CO(nC_st1_b182_c0));
  VFA U_st1_b182_c1 (.in_A(in_A[182]), .in_B(in_B[182]), .in_CI(1'b1), .out_S(nS_st1_b182_c1), .out_CO(nC_st1_b182_c1));
  VHA U_st1_b183_c0 (.in_A(in_A[183]), .in_B(in_B[183]), .out_S(nS_st1_b183_c0), .out_CO(nC_st1_b183_c0));
  VFA U_st1_b183_c1 (.in_A(in_A[183]), .in_B(in_B[183]), .in_CI(1'b1), .out_S(nS_st1_b183_c1), .out_CO(nC_st1_b183_c1));
  VHA U_st1_b184_c0 (.in_A(in_A[184]), .in_B(in_B[184]), .out_S(nS_st1_b184_c0), .out_CO(nC_st1_b184_c0));
  VFA U_st1_b184_c1 (.in_A(in_A[184]), .in_B(in_B[184]), .in_CI(1'b1), .out_S(nS_st1_b184_c1), .out_CO(nC_st1_b184_c1));
  VHA U_st1_b185_c0 (.in_A(in_A[185]), .in_B(in_B[185]), .out_S(nS_st1_b185_c0), .out_CO(nC_st1_b185_c0));
  VFA U_st1_b185_c1 (.in_A(in_A[185]), .in_B(in_B[185]), .in_CI(1'b1), .out_S(nS_st1_b185_c1), .out_CO(nC_st1_b185_c1));
  VHA U_st1_b186_c0 (.in_A(in_A[186]), .in_B(in_B[186]), .out_S(nS_st1_b186_c0), .out_CO(nC_st1_b186_c0));
  VFA U_st1_b186_c1 (.in_A(in_A[186]), .in_B(in_B[186]), .in_CI(1'b1), .out_S(nS_st1_b186_c1), .out_CO(nC_st1_b186_c1));
  VHA U_st1_b187_c0 (.in_A(in_A[187]), .in_B(in_B[187]), .out_S(nS_st1_b187_c0), .out_CO(nC_st1_b187_c0));
  VFA U_st1_b187_c1 (.in_A(in_A[187]), .in_B(in_B[187]), .in_CI(1'b1), .out_S(nS_st1_b187_c1), .out_CO(nC_st1_b187_c1));
  VHA U_st1_b188_c0 (.in_A(in_A[188]), .in_B(in_B[188]), .out_S(nS_st1_b188_c0), .out_CO(nC_st1_b188_c0));
  VFA U_st1_b188_c1 (.in_A(in_A[188]), .in_B(in_B[188]), .in_CI(1'b1), .out_S(nS_st1_b188_c1), .out_CO(nC_st1_b188_c1));
  VHA U_st1_b189_c0 (.in_A(in_A[189]), .in_B(in_B[189]), .out_S(nS_st1_b189_c0), .out_CO(nC_st1_b189_c0));
  VFA U_st1_b189_c1 (.in_A(in_A[189]), .in_B(in_B[189]), .in_CI(1'b1), .out_S(nS_st1_b189_c1), .out_CO(nC_st1_b189_c1));
  VHA U_st1_b190_c0 (.in_A(in_A[190]), .in_B(in_B[190]), .out_S(nS_st1_b190_c0), .out_CO(nC_st1_b190_c0));
  VFA U_st1_b190_c1 (.in_A(in_A[190]), .in_B(in_B[190]), .in_CI(1'b1), .out_S(nS_st1_b190_c1), .out_CO(nC_st1_b190_c1));
  VHA U_st1_b191_c0 (.in_A(in_A[191]), .in_B(in_B[191]), .out_S(nS_st1_b191_c0), .out_CO(nC_st1_b191_c0));
  VFA U_st1_b191_c1 (.in_A(in_A[191]), .in_B(in_B[191]), .in_CI(1'b1), .out_S(nS_st1_b191_c1), .out_CO(nC_st1_b191_c1));
  VHA U_st1_b192_c0 (.in_A(in_A[192]), .in_B(in_B[192]), .out_S(nS_st1_b192_c0), .out_CO(nC_st1_b192_c0));
  VFA U_st1_b192_c1 (.in_A(in_A[192]), .in_B(in_B[192]), .in_CI(1'b1), .out_S(nS_st1_b192_c1), .out_CO(nC_st1_b192_c1));
  VHA U_st1_b193_c0 (.in_A(in_A[193]), .in_B(in_B[193]), .out_S(nS_st1_b193_c0), .out_CO(nC_st1_b193_c0));
  VFA U_st1_b193_c1 (.in_A(in_A[193]), .in_B(in_B[193]), .in_CI(1'b1), .out_S(nS_st1_b193_c1), .out_CO(nC_st1_b193_c1));
  VHA U_st1_b194_c0 (.in_A(in_A[194]), .in_B(in_B[194]), .out_S(nS_st1_b194_c0), .out_CO(nC_st1_b194_c0));
  VFA U_st1_b194_c1 (.in_A(in_A[194]), .in_B(in_B[194]), .in_CI(1'b1), .out_S(nS_st1_b194_c1), .out_CO(nC_st1_b194_c1));
  VHA U_st1_b195_c0 (.in_A(in_A[195]), .in_B(in_B[195]), .out_S(nS_st1_b195_c0), .out_CO(nC_st1_b195_c0));
  VFA U_st1_b195_c1 (.in_A(in_A[195]), .in_B(in_B[195]), .in_CI(1'b1), .out_S(nS_st1_b195_c1), .out_CO(nC_st1_b195_c1));
  VHA U_st1_b196_c0 (.in_A(in_A[196]), .in_B(in_B[196]), .out_S(nS_st1_b196_c0), .out_CO(nC_st1_b196_c0));
  VFA U_st1_b196_c1 (.in_A(in_A[196]), .in_B(in_B[196]), .in_CI(1'b1), .out_S(nS_st1_b196_c1), .out_CO(nC_st1_b196_c1));
  VHA U_st1_b197_c0 (.in_A(in_A[197]), .in_B(in_B[197]), .out_S(nS_st1_b197_c0), .out_CO(nC_st1_b197_c0));
  VFA U_st1_b197_c1 (.in_A(in_A[197]), .in_B(in_B[197]), .in_CI(1'b1), .out_S(nS_st1_b197_c1), .out_CO(nC_st1_b197_c1));
  VHA U_st1_b198_c0 (.in_A(in_A[198]), .in_B(in_B[198]), .out_S(nS_st1_b198_c0), .out_CO(nC_st1_b198_c0));
  VFA U_st1_b198_c1 (.in_A(in_A[198]), .in_B(in_B[198]), .in_CI(1'b1), .out_S(nS_st1_b198_c1), .out_CO(nC_st1_b198_c1));
  VHA U_st1_b199_c0 (.in_A(in_A[199]), .in_B(in_B[199]), .out_S(nS_st1_b199_c0), .out_CO(nC_st1_b199_c0));
  VFA U_st1_b199_c1 (.in_A(in_A[199]), .in_B(in_B[199]), .in_CI(1'b1), .out_S(nS_st1_b199_c1), .out_CO(nC_st1_b199_c1));
  VHA U_st1_b200_c0 (.in_A(in_A[200]), .in_B(in_B[200]), .out_S(nS_st1_b200_c0), .out_CO(nC_st1_b200_c0));
  VFA U_st1_b200_c1 (.in_A(in_A[200]), .in_B(in_B[200]), .in_CI(1'b1), .out_S(nS_st1_b200_c1), .out_CO(nC_st1_b200_c1));
  VHA U_st1_b201_c0 (.in_A(in_A[201]), .in_B(in_B[201]), .out_S(nS_st1_b201_c0), .out_CO(nC_st1_b201_c0));
  VFA U_st1_b201_c1 (.in_A(in_A[201]), .in_B(in_B[201]), .in_CI(1'b1), .out_S(nS_st1_b201_c1), .out_CO(nC_st1_b201_c1));
  VHA U_st1_b202_c0 (.in_A(in_A[202]), .in_B(in_B[202]), .out_S(nS_st1_b202_c0), .out_CO(nC_st1_b202_c0));
  VFA U_st1_b202_c1 (.in_A(in_A[202]), .in_B(in_B[202]), .in_CI(1'b1), .out_S(nS_st1_b202_c1), .out_CO(nC_st1_b202_c1));
  VHA U_st1_b203_c0 (.in_A(in_A[203]), .in_B(in_B[203]), .out_S(nS_st1_b203_c0), .out_CO(nC_st1_b203_c0));
  VFA U_st1_b203_c1 (.in_A(in_A[203]), .in_B(in_B[203]), .in_CI(1'b1), .out_S(nS_st1_b203_c1), .out_CO(nC_st1_b203_c1));
  VHA U_st1_b204_c0 (.in_A(in_A[204]), .in_B(in_B[204]), .out_S(nS_st1_b204_c0), .out_CO(nC_st1_b204_c0));
  VFA U_st1_b204_c1 (.in_A(in_A[204]), .in_B(in_B[204]), .in_CI(1'b1), .out_S(nS_st1_b204_c1), .out_CO(nC_st1_b204_c1));
  VHA U_st1_b205_c0 (.in_A(in_A[205]), .in_B(in_B[205]), .out_S(nS_st1_b205_c0), .out_CO(nC_st1_b205_c0));
  VFA U_st1_b205_c1 (.in_A(in_A[205]), .in_B(in_B[205]), .in_CI(1'b1), .out_S(nS_st1_b205_c1), .out_CO(nC_st1_b205_c1));
  VHA U_st1_b206_c0 (.in_A(in_A[206]), .in_B(in_B[206]), .out_S(nS_st1_b206_c0), .out_CO(nC_st1_b206_c0));
  VFA U_st1_b206_c1 (.in_A(in_A[206]), .in_B(in_B[206]), .in_CI(1'b1), .out_S(nS_st1_b206_c1), .out_CO(nC_st1_b206_c1));
  VHA U_st1_b207_c0 (.in_A(in_A[207]), .in_B(in_B[207]), .out_S(nS_st1_b207_c0), .out_CO(nC_st1_b207_c0));
  VFA U_st1_b207_c1 (.in_A(in_A[207]), .in_B(in_B[207]), .in_CI(1'b1), .out_S(nS_st1_b207_c1), .out_CO(nC_st1_b207_c1));
  VHA U_st1_b208_c0 (.in_A(in_A[208]), .in_B(in_B[208]), .out_S(nS_st1_b208_c0), .out_CO(nC_st1_b208_c0));
  VFA U_st1_b208_c1 (.in_A(in_A[208]), .in_B(in_B[208]), .in_CI(1'b1), .out_S(nS_st1_b208_c1), .out_CO(nC_st1_b208_c1));
  VHA U_st1_b209_c0 (.in_A(in_A[209]), .in_B(in_B[209]), .out_S(nS_st1_b209_c0), .out_CO(nC_st1_b209_c0));
  VFA U_st1_b209_c1 (.in_A(in_A[209]), .in_B(in_B[209]), .in_CI(1'b1), .out_S(nS_st1_b209_c1), .out_CO(nC_st1_b209_c1));
  VHA U_st1_b210_c0 (.in_A(in_A[210]), .in_B(in_B[210]), .out_S(nS_st1_b210_c0), .out_CO(nC_st1_b210_c0));
  VFA U_st1_b210_c1 (.in_A(in_A[210]), .in_B(in_B[210]), .in_CI(1'b1), .out_S(nS_st1_b210_c1), .out_CO(nC_st1_b210_c1));
  VHA U_st1_b211_c0 (.in_A(in_A[211]), .in_B(in_B[211]), .out_S(nS_st1_b211_c0), .out_CO(nC_st1_b211_c0));
  VFA U_st1_b211_c1 (.in_A(in_A[211]), .in_B(in_B[211]), .in_CI(1'b1), .out_S(nS_st1_b211_c1), .out_CO(nC_st1_b211_c1));
  VHA U_st1_b212_c0 (.in_A(in_A[212]), .in_B(in_B[212]), .out_S(nS_st1_b212_c0), .out_CO(nC_st1_b212_c0));
  VFA U_st1_b212_c1 (.in_A(in_A[212]), .in_B(in_B[212]), .in_CI(1'b1), .out_S(nS_st1_b212_c1), .out_CO(nC_st1_b212_c1));
  VHA U_st1_b213_c0 (.in_A(in_A[213]), .in_B(in_B[213]), .out_S(nS_st1_b213_c0), .out_CO(nC_st1_b213_c0));
  VFA U_st1_b213_c1 (.in_A(in_A[213]), .in_B(in_B[213]), .in_CI(1'b1), .out_S(nS_st1_b213_c1), .out_CO(nC_st1_b213_c1));
  VHA U_st1_b214_c0 (.in_A(in_A[214]), .in_B(in_B[214]), .out_S(nS_st1_b214_c0), .out_CO(nC_st1_b214_c0));
  VFA U_st1_b214_c1 (.in_A(in_A[214]), .in_B(in_B[214]), .in_CI(1'b1), .out_S(nS_st1_b214_c1), .out_CO(nC_st1_b214_c1));
  VHA U_st1_b215_c0 (.in_A(in_A[215]), .in_B(in_B[215]), .out_S(nS_st1_b215_c0), .out_CO(nC_st1_b215_c0));
  VFA U_st1_b215_c1 (.in_A(in_A[215]), .in_B(in_B[215]), .in_CI(1'b1), .out_S(nS_st1_b215_c1), .out_CO(nC_st1_b215_c1));
  VHA U_st1_b216_c0 (.in_A(in_A[216]), .in_B(in_B[216]), .out_S(nS_st1_b216_c0), .out_CO(nC_st1_b216_c0));
  VFA U_st1_b216_c1 (.in_A(in_A[216]), .in_B(in_B[216]), .in_CI(1'b1), .out_S(nS_st1_b216_c1), .out_CO(nC_st1_b216_c1));
  VHA U_st1_b217_c0 (.in_A(in_A[217]), .in_B(in_B[217]), .out_S(nS_st1_b217_c0), .out_CO(nC_st1_b217_c0));
  VFA U_st1_b217_c1 (.in_A(in_A[217]), .in_B(in_B[217]), .in_CI(1'b1), .out_S(nS_st1_b217_c1), .out_CO(nC_st1_b217_c1));
  VHA U_st1_b218_c0 (.in_A(in_A[218]), .in_B(in_B[218]), .out_S(nS_st1_b218_c0), .out_CO(nC_st1_b218_c0));
  VFA U_st1_b218_c1 (.in_A(in_A[218]), .in_B(in_B[218]), .in_CI(1'b1), .out_S(nS_st1_b218_c1), .out_CO(nC_st1_b218_c1));
  VHA U_st1_b219_c0 (.in_A(in_A[219]), .in_B(in_B[219]), .out_S(nS_st1_b219_c0), .out_CO(nC_st1_b219_c0));
  VFA U_st1_b219_c1 (.in_A(in_A[219]), .in_B(in_B[219]), .in_CI(1'b1), .out_S(nS_st1_b219_c1), .out_CO(nC_st1_b219_c1));
  VHA U_st1_b220_c0 (.in_A(in_A[220]), .in_B(in_B[220]), .out_S(nS_st1_b220_c0), .out_CO(nC_st1_b220_c0));
  VFA U_st1_b220_c1 (.in_A(in_A[220]), .in_B(in_B[220]), .in_CI(1'b1), .out_S(nS_st1_b220_c1), .out_CO(nC_st1_b220_c1));
  VHA U_st1_b221_c0 (.in_A(in_A[221]), .in_B(in_B[221]), .out_S(nS_st1_b221_c0), .out_CO(nC_st1_b221_c0));
  VFA U_st1_b221_c1 (.in_A(in_A[221]), .in_B(in_B[221]), .in_CI(1'b1), .out_S(nS_st1_b221_c1), .out_CO(nC_st1_b221_c1));
  VHA U_st1_b222_c0 (.in_A(in_A[222]), .in_B(in_B[222]), .out_S(nS_st1_b222_c0), .out_CO(nC_st1_b222_c0));
  VFA U_st1_b222_c1 (.in_A(in_A[222]), .in_B(in_B[222]), .in_CI(1'b1), .out_S(nS_st1_b222_c1), .out_CO(nC_st1_b222_c1));
  VHA U_st1_b223_c0 (.in_A(in_A[223]), .in_B(in_B[223]), .out_S(nS_st1_b223_c0), .out_CO(nC_st1_b223_c0));
  VFA U_st1_b223_c1 (.in_A(in_A[223]), .in_B(in_B[223]), .in_CI(1'b1), .out_S(nS_st1_b223_c1), .out_CO(nC_st1_b223_c1));
  VHA U_st1_b224_c0 (.in_A(in_A[224]), .in_B(in_B[224]), .out_S(nS_st1_b224_c0), .out_CO(nC_st1_b224_c0));
  VFA U_st1_b224_c1 (.in_A(in_A[224]), .in_B(in_B[224]), .in_CI(1'b1), .out_S(nS_st1_b224_c1), .out_CO(nC_st1_b224_c1));
  VHA U_st1_b225_c0 (.in_A(in_A[225]), .in_B(in_B[225]), .out_S(nS_st1_b225_c0), .out_CO(nC_st1_b225_c0));
  VFA U_st1_b225_c1 (.in_A(in_A[225]), .in_B(in_B[225]), .in_CI(1'b1), .out_S(nS_st1_b225_c1), .out_CO(nC_st1_b225_c1));
  VHA U_st1_b226_c0 (.in_A(in_A[226]), .in_B(in_B[226]), .out_S(nS_st1_b226_c0), .out_CO(nC_st1_b226_c0));
  VFA U_st1_b226_c1 (.in_A(in_A[226]), .in_B(in_B[226]), .in_CI(1'b1), .out_S(nS_st1_b226_c1), .out_CO(nC_st1_b226_c1));
  VHA U_st1_b227_c0 (.in_A(in_A[227]), .in_B(in_B[227]), .out_S(nS_st1_b227_c0), .out_CO(nC_st1_b227_c0));
  VFA U_st1_b227_c1 (.in_A(in_A[227]), .in_B(in_B[227]), .in_CI(1'b1), .out_S(nS_st1_b227_c1), .out_CO(nC_st1_b227_c1));
  VHA U_st1_b228_c0 (.in_A(in_A[228]), .in_B(in_B[228]), .out_S(nS_st1_b228_c0), .out_CO(nC_st1_b228_c0));
  VFA U_st1_b228_c1 (.in_A(in_A[228]), .in_B(in_B[228]), .in_CI(1'b1), .out_S(nS_st1_b228_c1), .out_CO(nC_st1_b228_c1));
  VHA U_st1_b229_c0 (.in_A(in_A[229]), .in_B(in_B[229]), .out_S(nS_st1_b229_c0), .out_CO(nC_st1_b229_c0));
  VFA U_st1_b229_c1 (.in_A(in_A[229]), .in_B(in_B[229]), .in_CI(1'b1), .out_S(nS_st1_b229_c1), .out_CO(nC_st1_b229_c1));
  VHA U_st1_b230_c0 (.in_A(in_A[230]), .in_B(in_B[230]), .out_S(nS_st1_b230_c0), .out_CO(nC_st1_b230_c0));
  VFA U_st1_b230_c1 (.in_A(in_A[230]), .in_B(in_B[230]), .in_CI(1'b1), .out_S(nS_st1_b230_c1), .out_CO(nC_st1_b230_c1));
  VHA U_st1_b231_c0 (.in_A(in_A[231]), .in_B(in_B[231]), .out_S(nS_st1_b231_c0), .out_CO(nC_st1_b231_c0));
  VFA U_st1_b231_c1 (.in_A(in_A[231]), .in_B(in_B[231]), .in_CI(1'b1), .out_S(nS_st1_b231_c1), .out_CO(nC_st1_b231_c1));
  VHA U_st1_b232_c0 (.in_A(in_A[232]), .in_B(in_B[232]), .out_S(nS_st1_b232_c0), .out_CO(nC_st1_b232_c0));
  VFA U_st1_b232_c1 (.in_A(in_A[232]), .in_B(in_B[232]), .in_CI(1'b1), .out_S(nS_st1_b232_c1), .out_CO(nC_st1_b232_c1));
  VHA U_st1_b233_c0 (.in_A(in_A[233]), .in_B(in_B[233]), .out_S(nS_st1_b233_c0), .out_CO(nC_st1_b233_c0));
  VFA U_st1_b233_c1 (.in_A(in_A[233]), .in_B(in_B[233]), .in_CI(1'b1), .out_S(nS_st1_b233_c1), .out_CO(nC_st1_b233_c1));
  VHA U_st1_b234_c0 (.in_A(in_A[234]), .in_B(in_B[234]), .out_S(nS_st1_b234_c0), .out_CO(nC_st1_b234_c0));
  VFA U_st1_b234_c1 (.in_A(in_A[234]), .in_B(in_B[234]), .in_CI(1'b1), .out_S(nS_st1_b234_c1), .out_CO(nC_st1_b234_c1));
  VHA U_st1_b235_c0 (.in_A(in_A[235]), .in_B(in_B[235]), .out_S(nS_st1_b235_c0), .out_CO(nC_st1_b235_c0));
  VFA U_st1_b235_c1 (.in_A(in_A[235]), .in_B(in_B[235]), .in_CI(1'b1), .out_S(nS_st1_b235_c1), .out_CO(nC_st1_b235_c1));
  VHA U_st1_b236_c0 (.in_A(in_A[236]), .in_B(in_B[236]), .out_S(nS_st1_b236_c0), .out_CO(nC_st1_b236_c0));
  VFA U_st1_b236_c1 (.in_A(in_A[236]), .in_B(in_B[236]), .in_CI(1'b1), .out_S(nS_st1_b236_c1), .out_CO(nC_st1_b236_c1));
  VHA U_st1_b237_c0 (.in_A(in_A[237]), .in_B(in_B[237]), .out_S(nS_st1_b237_c0), .out_CO(nC_st1_b237_c0));
  VFA U_st1_b237_c1 (.in_A(in_A[237]), .in_B(in_B[237]), .in_CI(1'b1), .out_S(nS_st1_b237_c1), .out_CO(nC_st1_b237_c1));
  VHA U_st1_b238_c0 (.in_A(in_A[238]), .in_B(in_B[238]), .out_S(nS_st1_b238_c0), .out_CO(nC_st1_b238_c0));
  VFA U_st1_b238_c1 (.in_A(in_A[238]), .in_B(in_B[238]), .in_CI(1'b1), .out_S(nS_st1_b238_c1), .out_CO(nC_st1_b238_c1));
  VHA U_st1_b239_c0 (.in_A(in_A[239]), .in_B(in_B[239]), .out_S(nS_st1_b239_c0), .out_CO(nC_st1_b239_c0));
  VFA U_st1_b239_c1 (.in_A(in_A[239]), .in_B(in_B[239]), .in_CI(1'b1), .out_S(nS_st1_b239_c1), .out_CO(nC_st1_b239_c1));
  VHA U_st1_b240_c0 (.in_A(in_A[240]), .in_B(in_B[240]), .out_S(nS_st1_b240_c0), .out_CO(nC_st1_b240_c0));
  VFA U_st1_b240_c1 (.in_A(in_A[240]), .in_B(in_B[240]), .in_CI(1'b1), .out_S(nS_st1_b240_c1), .out_CO(nC_st1_b240_c1));
  VHA U_st1_b241_c0 (.in_A(in_A[241]), .in_B(in_B[241]), .out_S(nS_st1_b241_c0), .out_CO(nC_st1_b241_c0));
  VFA U_st1_b241_c1 (.in_A(in_A[241]), .in_B(in_B[241]), .in_CI(1'b1), .out_S(nS_st1_b241_c1), .out_CO(nC_st1_b241_c1));
  VHA U_st1_b242_c0 (.in_A(in_A[242]), .in_B(in_B[242]), .out_S(nS_st1_b242_c0), .out_CO(nC_st1_b242_c0));
  VFA U_st1_b242_c1 (.in_A(in_A[242]), .in_B(in_B[242]), .in_CI(1'b1), .out_S(nS_st1_b242_c1), .out_CO(nC_st1_b242_c1));
  VHA U_st1_b243_c0 (.in_A(in_A[243]), .in_B(in_B[243]), .out_S(nS_st1_b243_c0), .out_CO(nC_st1_b243_c0));
  VFA U_st1_b243_c1 (.in_A(in_A[243]), .in_B(in_B[243]), .in_CI(1'b1), .out_S(nS_st1_b243_c1), .out_CO(nC_st1_b243_c1));
  VHA U_st1_b244_c0 (.in_A(in_A[244]), .in_B(in_B[244]), .out_S(nS_st1_b244_c0), .out_CO(nC_st1_b244_c0));
  VFA U_st1_b244_c1 (.in_A(in_A[244]), .in_B(in_B[244]), .in_CI(1'b1), .out_S(nS_st1_b244_c1), .out_CO(nC_st1_b244_c1));
  VHA U_st1_b245_c0 (.in_A(in_A[245]), .in_B(in_B[245]), .out_S(nS_st1_b245_c0), .out_CO(nC_st1_b245_c0));
  VFA U_st1_b245_c1 (.in_A(in_A[245]), .in_B(in_B[245]), .in_CI(1'b1), .out_S(nS_st1_b245_c1), .out_CO(nC_st1_b245_c1));
  VHA U_st1_b246_c0 (.in_A(in_A[246]), .in_B(in_B[246]), .out_S(nS_st1_b246_c0), .out_CO(nC_st1_b246_c0));
  VFA U_st1_b246_c1 (.in_A(in_A[246]), .in_B(in_B[246]), .in_CI(1'b1), .out_S(nS_st1_b246_c1), .out_CO(nC_st1_b246_c1));
  VHA U_st1_b247_c0 (.in_A(in_A[247]), .in_B(in_B[247]), .out_S(nS_st1_b247_c0), .out_CO(nC_st1_b247_c0));
  VFA U_st1_b247_c1 (.in_A(in_A[247]), .in_B(in_B[247]), .in_CI(1'b1), .out_S(nS_st1_b247_c1), .out_CO(nC_st1_b247_c1));
  VHA U_st1_b248_c0 (.in_A(in_A[248]), .in_B(in_B[248]), .out_S(nS_st1_b248_c0), .out_CO(nC_st1_b248_c0));
  VFA U_st1_b248_c1 (.in_A(in_A[248]), .in_B(in_B[248]), .in_CI(1'b1), .out_S(nS_st1_b248_c1), .out_CO(nC_st1_b248_c1));
  VHA U_st1_b249_c0 (.in_A(in_A[249]), .in_B(in_B[249]), .out_S(nS_st1_b249_c0), .out_CO(nC_st1_b249_c0));
  VFA U_st1_b249_c1 (.in_A(in_A[249]), .in_B(in_B[249]), .in_CI(1'b1), .out_S(nS_st1_b249_c1), .out_CO(nC_st1_b249_c1));
  VHA U_st1_b250_c0 (.in_A(in_A[250]), .in_B(in_B[250]), .out_S(nS_st1_b250_c0), .out_CO(nC_st1_b250_c0));
  VFA U_st1_b250_c1 (.in_A(in_A[250]), .in_B(in_B[250]), .in_CI(1'b1), .out_S(nS_st1_b250_c1), .out_CO(nC_st1_b250_c1));
  VHA U_st1_b251_c0 (.in_A(in_A[251]), .in_B(in_B[251]), .out_S(nS_st1_b251_c0), .out_CO(nC_st1_b251_c0));
  VFA U_st1_b251_c1 (.in_A(in_A[251]), .in_B(in_B[251]), .in_CI(1'b1), .out_S(nS_st1_b251_c1), .out_CO(nC_st1_b251_c1));
  VHA U_st1_b252_c0 (.in_A(in_A[252]), .in_B(in_B[252]), .out_S(nS_st1_b252_c0), .out_CO(nC_st1_b252_c0));
  VFA U_st1_b252_c1 (.in_A(in_A[252]), .in_B(in_B[252]), .in_CI(1'b1), .out_S(nS_st1_b252_c1), .out_CO(nC_st1_b252_c1));
  VHA U_st1_b253_c0 (.in_A(in_A[253]), .in_B(in_B[253]), .out_S(nS_st1_b253_c0), .out_CO(nC_st1_b253_c0));
  VFA U_st1_b253_c1 (.in_A(in_A[253]), .in_B(in_B[253]), .in_CI(1'b1), .out_S(nS_st1_b253_c1), .out_CO(nC_st1_b253_c1));
  VHA U_st1_b254_c0 (.in_A(in_A[254]), .in_B(in_B[254]), .out_S(nS_st1_b254_c0), .out_CO(nC_st1_b254_c0));
  VFA U_st1_b254_c1 (.in_A(in_A[254]), .in_B(in_B[254]), .in_CI(1'b1), .out_S(nS_st1_b254_c1), .out_CO(nC_st1_b254_c1));
  VHA U_st1_b255_c0 (.in_A(in_A[255]), .in_B(in_B[255]), .out_S(nS_st1_b255_c0), .out_CO(nC_st1_b255_c0));
  VFA U_st1_b255_c1 (.in_A(in_A[255]), .in_B(in_B[255]), .in_CI(1'b1), .out_S(nS_st1_b255_c1), .out_CO(nC_st1_b255_c1));

  assign nS_st2_b0_c0 = nS_st1_b0_c0;
  assign nS_st2_b1_c0 = (nC_st1_b0_c0 == 0) ? nS_st1_b1_c0 : nS_st1_b1_c1;
  assign nS_st2_b2_c0 = nS_st1_b2_c0;
  assign nS_st2_b3_c0 = (nC_st1_b2_c0 == 0) ? nS_st1_b3_c0 : nS_st1_b3_c1;
  assign nS_st2_b4_c0 = nS_st1_b4_c0;
  assign nS_st2_b5_c0 = (nC_st1_b4_c0 == 0) ? nS_st1_b5_c0 : nS_st1_b5_c1;
  assign nS_st2_b6_c0 = nS_st1_b6_c0;
  assign nS_st2_b7_c0 = (nC_st1_b6_c0 == 0) ? nS_st1_b7_c0 : nS_st1_b7_c1;
  assign nS_st2_b8_c0 = nS_st1_b8_c0;
  assign nS_st2_b9_c0 = (nC_st1_b8_c0 == 0) ? nS_st1_b9_c0 : nS_st1_b9_c1;
  assign nS_st2_b10_c0 = nS_st1_b10_c0;
  assign nS_st2_b11_c0 = (nC_st1_b10_c0 == 0) ? nS_st1_b11_c0 : nS_st1_b11_c1;
  assign nS_st2_b12_c0 = nS_st1_b12_c0;
  assign nS_st2_b13_c0 = (nC_st1_b12_c0 == 0) ? nS_st1_b13_c0 : nS_st1_b13_c1;
  assign nS_st2_b14_c0 = nS_st1_b14_c0;
  assign nS_st2_b15_c0 = (nC_st1_b14_c0 == 0) ? nS_st1_b15_c0 : nS_st1_b15_c1;
  assign nS_st2_b16_c0 = nS_st1_b16_c0;
  assign nS_st2_b17_c0 = (nC_st1_b16_c0 == 0) ? nS_st1_b17_c0 : nS_st1_b17_c1;
  assign nS_st2_b18_c0 = nS_st1_b18_c0;
  assign nS_st2_b19_c0 = (nC_st1_b18_c0 == 0) ? nS_st1_b19_c0 : nS_st1_b19_c1;
  assign nS_st2_b20_c0 = nS_st1_b20_c0;
  assign nS_st2_b21_c0 = (nC_st1_b20_c0 == 0) ? nS_st1_b21_c0 : nS_st1_b21_c1;
  assign nS_st2_b22_c0 = nS_st1_b22_c0;
  assign nS_st2_b23_c0 = (nC_st1_b22_c0 == 0) ? nS_st1_b23_c0 : nS_st1_b23_c1;
  assign nS_st2_b24_c0 = nS_st1_b24_c0;
  assign nS_st2_b25_c0 = (nC_st1_b24_c0 == 0) ? nS_st1_b25_c0 : nS_st1_b25_c1;
  assign nS_st2_b26_c0 = nS_st1_b26_c0;
  assign nS_st2_b27_c0 = (nC_st1_b26_c0 == 0) ? nS_st1_b27_c0 : nS_st1_b27_c1;
  assign nS_st2_b28_c0 = nS_st1_b28_c0;
  assign nS_st2_b29_c0 = (nC_st1_b28_c0 == 0) ? nS_st1_b29_c0 : nS_st1_b29_c1;
  assign nS_st2_b30_c0 = nS_st1_b30_c0;
  assign nS_st2_b31_c0 = (nC_st1_b30_c0 == 0) ? nS_st1_b31_c0 : nS_st1_b31_c1;
  assign nS_st2_b32_c0 = nS_st1_b32_c0;
  assign nS_st2_b33_c0 = (nC_st1_b32_c0 == 0) ? nS_st1_b33_c0 : nS_st1_b33_c1;
  assign nS_st2_b34_c0 = nS_st1_b34_c0;
  assign nS_st2_b35_c0 = (nC_st1_b34_c0 == 0) ? nS_st1_b35_c0 : nS_st1_b35_c1;
  assign nS_st2_b36_c0 = nS_st1_b36_c0;
  assign nS_st2_b37_c0 = (nC_st1_b36_c0 == 0) ? nS_st1_b37_c0 : nS_st1_b37_c1;
  assign nS_st2_b38_c0 = nS_st1_b38_c0;
  assign nS_st2_b39_c0 = (nC_st1_b38_c0 == 0) ? nS_st1_b39_c0 : nS_st1_b39_c1;
  assign nS_st2_b40_c0 = nS_st1_b40_c0;
  assign nS_st2_b41_c0 = (nC_st1_b40_c0 == 0) ? nS_st1_b41_c0 : nS_st1_b41_c1;
  assign nS_st2_b42_c0 = nS_st1_b42_c0;
  assign nS_st2_b43_c0 = (nC_st1_b42_c0 == 0) ? nS_st1_b43_c0 : nS_st1_b43_c1;
  assign nS_st2_b44_c0 = nS_st1_b44_c0;
  assign nS_st2_b45_c0 = (nC_st1_b44_c0 == 0) ? nS_st1_b45_c0 : nS_st1_b45_c1;
  assign nS_st2_b46_c0 = nS_st1_b46_c0;
  assign nS_st2_b47_c0 = (nC_st1_b46_c0 == 0) ? nS_st1_b47_c0 : nS_st1_b47_c1;
  assign nS_st2_b48_c0 = nS_st1_b48_c0;
  assign nS_st2_b49_c0 = (nC_st1_b48_c0 == 0) ? nS_st1_b49_c0 : nS_st1_b49_c1;
  assign nS_st2_b50_c0 = nS_st1_b50_c0;
  assign nS_st2_b51_c0 = (nC_st1_b50_c0 == 0) ? nS_st1_b51_c0 : nS_st1_b51_c1;
  assign nS_st2_b52_c0 = nS_st1_b52_c0;
  assign nS_st2_b53_c0 = (nC_st1_b52_c0 == 0) ? nS_st1_b53_c0 : nS_st1_b53_c1;
  assign nS_st2_b54_c0 = nS_st1_b54_c0;
  assign nS_st2_b55_c0 = (nC_st1_b54_c0 == 0) ? nS_st1_b55_c0 : nS_st1_b55_c1;
  assign nS_st2_b56_c0 = nS_st1_b56_c0;
  assign nS_st2_b57_c0 = (nC_st1_b56_c0 == 0) ? nS_st1_b57_c0 : nS_st1_b57_c1;
  assign nS_st2_b58_c0 = nS_st1_b58_c0;
  assign nS_st2_b59_c0 = (nC_st1_b58_c0 == 0) ? nS_st1_b59_c0 : nS_st1_b59_c1;
  assign nS_st2_b60_c0 = nS_st1_b60_c0;
  assign nS_st2_b61_c0 = (nC_st1_b60_c0 == 0) ? nS_st1_b61_c0 : nS_st1_b61_c1;
  assign nS_st2_b62_c0 = nS_st1_b62_c0;
  assign nS_st2_b63_c0 = (nC_st1_b62_c0 == 0) ? nS_st1_b63_c0 : nS_st1_b63_c1;
  assign nS_st2_b64_c0 = nS_st1_b64_c0;
  assign nS_st2_b65_c0 = (nC_st1_b64_c0 == 0) ? nS_st1_b65_c0 : nS_st1_b65_c1;
  assign nS_st2_b66_c0 = nS_st1_b66_c0;
  assign nS_st2_b67_c0 = (nC_st1_b66_c0 == 0) ? nS_st1_b67_c0 : nS_st1_b67_c1;
  assign nS_st2_b68_c0 = nS_st1_b68_c0;
  assign nS_st2_b69_c0 = (nC_st1_b68_c0 == 0) ? nS_st1_b69_c0 : nS_st1_b69_c1;
  assign nS_st2_b70_c0 = nS_st1_b70_c0;
  assign nS_st2_b71_c0 = (nC_st1_b70_c0 == 0) ? nS_st1_b71_c0 : nS_st1_b71_c1;
  assign nS_st2_b72_c0 = nS_st1_b72_c0;
  assign nS_st2_b73_c0 = (nC_st1_b72_c0 == 0) ? nS_st1_b73_c0 : nS_st1_b73_c1;
  assign nS_st2_b74_c0 = nS_st1_b74_c0;
  assign nS_st2_b75_c0 = (nC_st1_b74_c0 == 0) ? nS_st1_b75_c0 : nS_st1_b75_c1;
  assign nS_st2_b76_c0 = nS_st1_b76_c0;
  assign nS_st2_b77_c0 = (nC_st1_b76_c0 == 0) ? nS_st1_b77_c0 : nS_st1_b77_c1;
  assign nS_st2_b78_c0 = nS_st1_b78_c0;
  assign nS_st2_b79_c0 = (nC_st1_b78_c0 == 0) ? nS_st1_b79_c0 : nS_st1_b79_c1;
  assign nS_st2_b80_c0 = nS_st1_b80_c0;
  assign nS_st2_b81_c0 = (nC_st1_b80_c0 == 0) ? nS_st1_b81_c0 : nS_st1_b81_c1;
  assign nS_st2_b82_c0 = nS_st1_b82_c0;
  assign nS_st2_b83_c0 = (nC_st1_b82_c0 == 0) ? nS_st1_b83_c0 : nS_st1_b83_c1;
  assign nS_st2_b84_c0 = nS_st1_b84_c0;
  assign nS_st2_b85_c0 = (nC_st1_b84_c0 == 0) ? nS_st1_b85_c0 : nS_st1_b85_c1;
  assign nS_st2_b86_c0 = nS_st1_b86_c0;
  assign nS_st2_b87_c0 = (nC_st1_b86_c0 == 0) ? nS_st1_b87_c0 : nS_st1_b87_c1;
  assign nS_st2_b88_c0 = nS_st1_b88_c0;
  assign nS_st2_b89_c0 = (nC_st1_b88_c0 == 0) ? nS_st1_b89_c0 : nS_st1_b89_c1;
  assign nS_st2_b90_c0 = nS_st1_b90_c0;
  assign nS_st2_b91_c0 = (nC_st1_b90_c0 == 0) ? nS_st1_b91_c0 : nS_st1_b91_c1;
  assign nS_st2_b92_c0 = nS_st1_b92_c0;
  assign nS_st2_b93_c0 = (nC_st1_b92_c0 == 0) ? nS_st1_b93_c0 : nS_st1_b93_c1;
  assign nS_st2_b94_c0 = nS_st1_b94_c0;
  assign nS_st2_b95_c0 = (nC_st1_b94_c0 == 0) ? nS_st1_b95_c0 : nS_st1_b95_c1;
  assign nS_st2_b96_c0 = nS_st1_b96_c0;
  assign nS_st2_b97_c0 = (nC_st1_b96_c0 == 0) ? nS_st1_b97_c0 : nS_st1_b97_c1;
  assign nS_st2_b98_c0 = nS_st1_b98_c0;
  assign nS_st2_b99_c0 = (nC_st1_b98_c0 == 0) ? nS_st1_b99_c0 : nS_st1_b99_c1;
  assign nS_st2_b100_c0 = nS_st1_b100_c0;
  assign nS_st2_b101_c0 = (nC_st1_b100_c0 == 0) ? nS_st1_b101_c0 : nS_st1_b101_c1;
  assign nS_st2_b102_c0 = nS_st1_b102_c0;
  assign nS_st2_b103_c0 = (nC_st1_b102_c0 == 0) ? nS_st1_b103_c0 : nS_st1_b103_c1;
  assign nS_st2_b104_c0 = nS_st1_b104_c0;
  assign nS_st2_b105_c0 = (nC_st1_b104_c0 == 0) ? nS_st1_b105_c0 : nS_st1_b105_c1;
  assign nS_st2_b106_c0 = nS_st1_b106_c0;
  assign nS_st2_b107_c0 = (nC_st1_b106_c0 == 0) ? nS_st1_b107_c0 : nS_st1_b107_c1;
  assign nS_st2_b108_c0 = nS_st1_b108_c0;
  assign nS_st2_b109_c0 = (nC_st1_b108_c0 == 0) ? nS_st1_b109_c0 : nS_st1_b109_c1;
  assign nS_st2_b110_c0 = nS_st1_b110_c0;
  assign nS_st2_b111_c0 = (nC_st1_b110_c0 == 0) ? nS_st1_b111_c0 : nS_st1_b111_c1;
  assign nS_st2_b112_c0 = nS_st1_b112_c0;
  assign nS_st2_b113_c0 = (nC_st1_b112_c0 == 0) ? nS_st1_b113_c0 : nS_st1_b113_c1;
  assign nS_st2_b114_c0 = nS_st1_b114_c0;
  assign nS_st2_b115_c0 = (nC_st1_b114_c0 == 0) ? nS_st1_b115_c0 : nS_st1_b115_c1;
  assign nS_st2_b116_c0 = nS_st1_b116_c0;
  assign nS_st2_b117_c0 = (nC_st1_b116_c0 == 0) ? nS_st1_b117_c0 : nS_st1_b117_c1;
  assign nS_st2_b118_c0 = nS_st1_b118_c0;
  assign nS_st2_b119_c0 = (nC_st1_b118_c0 == 0) ? nS_st1_b119_c0 : nS_st1_b119_c1;
  assign nS_st2_b120_c0 = nS_st1_b120_c0;
  assign nS_st2_b121_c0 = (nC_st1_b120_c0 == 0) ? nS_st1_b121_c0 : nS_st1_b121_c1;
  assign nS_st2_b122_c0 = nS_st1_b122_c0;
  assign nS_st2_b123_c0 = (nC_st1_b122_c0 == 0) ? nS_st1_b123_c0 : nS_st1_b123_c1;
  assign nS_st2_b124_c0 = nS_st1_b124_c0;
  assign nS_st2_b125_c0 = (nC_st1_b124_c0 == 0) ? nS_st1_b125_c0 : nS_st1_b125_c1;
  assign nS_st2_b126_c0 = nS_st1_b126_c0;
  assign nS_st2_b127_c0 = (nC_st1_b126_c0 == 0) ? nS_st1_b127_c0 : nS_st1_b127_c1;
  assign nS_st2_b128_c0 = nS_st1_b128_c0;
  assign nS_st2_b129_c0 = (nC_st1_b128_c0 == 0) ? nS_st1_b129_c0 : nS_st1_b129_c1;
  assign nS_st2_b130_c0 = nS_st1_b130_c0;
  assign nS_st2_b131_c0 = (nC_st1_b130_c0 == 0) ? nS_st1_b131_c0 : nS_st1_b131_c1;
  assign nS_st2_b132_c0 = nS_st1_b132_c0;
  assign nS_st2_b133_c0 = (nC_st1_b132_c0 == 0) ? nS_st1_b133_c0 : nS_st1_b133_c1;
  assign nS_st2_b134_c0 = nS_st1_b134_c0;
  assign nS_st2_b135_c0 = (nC_st1_b134_c0 == 0) ? nS_st1_b135_c0 : nS_st1_b135_c1;
  assign nS_st2_b136_c0 = nS_st1_b136_c0;
  assign nS_st2_b137_c0 = (nC_st1_b136_c0 == 0) ? nS_st1_b137_c0 : nS_st1_b137_c1;
  assign nS_st2_b138_c0 = nS_st1_b138_c0;
  assign nS_st2_b139_c0 = (nC_st1_b138_c0 == 0) ? nS_st1_b139_c0 : nS_st1_b139_c1;
  assign nS_st2_b140_c0 = nS_st1_b140_c0;
  assign nS_st2_b141_c0 = (nC_st1_b140_c0 == 0) ? nS_st1_b141_c0 : nS_st1_b141_c1;
  assign nS_st2_b142_c0 = nS_st1_b142_c0;
  assign nS_st2_b143_c0 = (nC_st1_b142_c0 == 0) ? nS_st1_b143_c0 : nS_st1_b143_c1;
  assign nS_st2_b144_c0 = nS_st1_b144_c0;
  assign nS_st2_b145_c0 = (nC_st1_b144_c0 == 0) ? nS_st1_b145_c0 : nS_st1_b145_c1;
  assign nS_st2_b146_c0 = nS_st1_b146_c0;
  assign nS_st2_b147_c0 = (nC_st1_b146_c0 == 0) ? nS_st1_b147_c0 : nS_st1_b147_c1;
  assign nS_st2_b148_c0 = nS_st1_b148_c0;
  assign nS_st2_b149_c0 = (nC_st1_b148_c0 == 0) ? nS_st1_b149_c0 : nS_st1_b149_c1;
  assign nS_st2_b150_c0 = nS_st1_b150_c0;
  assign nS_st2_b151_c0 = (nC_st1_b150_c0 == 0) ? nS_st1_b151_c0 : nS_st1_b151_c1;
  assign nS_st2_b152_c0 = nS_st1_b152_c0;
  assign nS_st2_b153_c0 = (nC_st1_b152_c0 == 0) ? nS_st1_b153_c0 : nS_st1_b153_c1;
  assign nS_st2_b154_c0 = nS_st1_b154_c0;
  assign nS_st2_b155_c0 = (nC_st1_b154_c0 == 0) ? nS_st1_b155_c0 : nS_st1_b155_c1;
  assign nS_st2_b156_c0 = nS_st1_b156_c0;
  assign nS_st2_b157_c0 = (nC_st1_b156_c0 == 0) ? nS_st1_b157_c0 : nS_st1_b157_c1;
  assign nS_st2_b158_c0 = nS_st1_b158_c0;
  assign nS_st2_b159_c0 = (nC_st1_b158_c0 == 0) ? nS_st1_b159_c0 : nS_st1_b159_c1;
  assign nS_st2_b160_c0 = nS_st1_b160_c0;
  assign nS_st2_b161_c0 = (nC_st1_b160_c0 == 0) ? nS_st1_b161_c0 : nS_st1_b161_c1;
  assign nS_st2_b162_c0 = nS_st1_b162_c0;
  assign nS_st2_b163_c0 = (nC_st1_b162_c0 == 0) ? nS_st1_b163_c0 : nS_st1_b163_c1;
  assign nS_st2_b164_c0 = nS_st1_b164_c0;
  assign nS_st2_b165_c0 = (nC_st1_b164_c0 == 0) ? nS_st1_b165_c0 : nS_st1_b165_c1;
  assign nS_st2_b166_c0 = nS_st1_b166_c0;
  assign nS_st2_b167_c0 = (nC_st1_b166_c0 == 0) ? nS_st1_b167_c0 : nS_st1_b167_c1;
  assign nS_st2_b168_c0 = nS_st1_b168_c0;
  assign nS_st2_b169_c0 = (nC_st1_b168_c0 == 0) ? nS_st1_b169_c0 : nS_st1_b169_c1;
  assign nS_st2_b170_c0 = nS_st1_b170_c0;
  assign nS_st2_b171_c0 = (nC_st1_b170_c0 == 0) ? nS_st1_b171_c0 : nS_st1_b171_c1;
  assign nS_st2_b172_c0 = nS_st1_b172_c0;
  assign nS_st2_b173_c0 = (nC_st1_b172_c0 == 0) ? nS_st1_b173_c0 : nS_st1_b173_c1;
  assign nS_st2_b174_c0 = nS_st1_b174_c0;
  assign nS_st2_b175_c0 = (nC_st1_b174_c0 == 0) ? nS_st1_b175_c0 : nS_st1_b175_c1;
  assign nS_st2_b176_c0 = nS_st1_b176_c0;
  assign nS_st2_b177_c0 = (nC_st1_b176_c0 == 0) ? nS_st1_b177_c0 : nS_st1_b177_c1;
  assign nS_st2_b178_c0 = nS_st1_b178_c0;
  assign nS_st2_b179_c0 = (nC_st1_b178_c0 == 0) ? nS_st1_b179_c0 : nS_st1_b179_c1;
  assign nS_st2_b180_c0 = nS_st1_b180_c0;
  assign nS_st2_b181_c0 = (nC_st1_b180_c0 == 0) ? nS_st1_b181_c0 : nS_st1_b181_c1;
  assign nS_st2_b182_c0 = nS_st1_b182_c0;
  assign nS_st2_b183_c0 = (nC_st1_b182_c0 == 0) ? nS_st1_b183_c0 : nS_st1_b183_c1;
  assign nS_st2_b184_c0 = nS_st1_b184_c0;
  assign nS_st2_b185_c0 = (nC_st1_b184_c0 == 0) ? nS_st1_b185_c0 : nS_st1_b185_c1;
  assign nS_st2_b186_c0 = nS_st1_b186_c0;
  assign nS_st2_b187_c0 = (nC_st1_b186_c0 == 0) ? nS_st1_b187_c0 : nS_st1_b187_c1;
  assign nS_st2_b188_c0 = nS_st1_b188_c0;
  assign nS_st2_b189_c0 = (nC_st1_b188_c0 == 0) ? nS_st1_b189_c0 : nS_st1_b189_c1;
  assign nS_st2_b190_c0 = nS_st1_b190_c0;
  assign nS_st2_b191_c0 = (nC_st1_b190_c0 == 0) ? nS_st1_b191_c0 : nS_st1_b191_c1;
  assign nS_st2_b192_c0 = nS_st1_b192_c0;
  assign nS_st2_b193_c0 = (nC_st1_b192_c0 == 0) ? nS_st1_b193_c0 : nS_st1_b193_c1;
  assign nS_st2_b194_c0 = nS_st1_b194_c0;
  assign nS_st2_b195_c0 = (nC_st1_b194_c0 == 0) ? nS_st1_b195_c0 : nS_st1_b195_c1;
  assign nS_st2_b196_c0 = nS_st1_b196_c0;
  assign nS_st2_b197_c0 = (nC_st1_b196_c0 == 0) ? nS_st1_b197_c0 : nS_st1_b197_c1;
  assign nS_st2_b198_c0 = nS_st1_b198_c0;
  assign nS_st2_b199_c0 = (nC_st1_b198_c0 == 0) ? nS_st1_b199_c0 : nS_st1_b199_c1;
  assign nS_st2_b200_c0 = nS_st1_b200_c0;
  assign nS_st2_b201_c0 = (nC_st1_b200_c0 == 0) ? nS_st1_b201_c0 : nS_st1_b201_c1;
  assign nS_st2_b202_c0 = nS_st1_b202_c0;
  assign nS_st2_b203_c0 = (nC_st1_b202_c0 == 0) ? nS_st1_b203_c0 : nS_st1_b203_c1;
  assign nS_st2_b204_c0 = nS_st1_b204_c0;
  assign nS_st2_b205_c0 = (nC_st1_b204_c0 == 0) ? nS_st1_b205_c0 : nS_st1_b205_c1;
  assign nS_st2_b206_c0 = nS_st1_b206_c0;
  assign nS_st2_b207_c0 = (nC_st1_b206_c0 == 0) ? nS_st1_b207_c0 : nS_st1_b207_c1;
  assign nS_st2_b208_c0 = nS_st1_b208_c0;
  assign nS_st2_b209_c0 = (nC_st1_b208_c0 == 0) ? nS_st1_b209_c0 : nS_st1_b209_c1;
  assign nS_st2_b210_c0 = nS_st1_b210_c0;
  assign nS_st2_b211_c0 = (nC_st1_b210_c0 == 0) ? nS_st1_b211_c0 : nS_st1_b211_c1;
  assign nS_st2_b212_c0 = nS_st1_b212_c0;
  assign nS_st2_b213_c0 = (nC_st1_b212_c0 == 0) ? nS_st1_b213_c0 : nS_st1_b213_c1;
  assign nS_st2_b214_c0 = nS_st1_b214_c0;
  assign nS_st2_b215_c0 = (nC_st1_b214_c0 == 0) ? nS_st1_b215_c0 : nS_st1_b215_c1;
  assign nS_st2_b216_c0 = nS_st1_b216_c0;
  assign nS_st2_b217_c0 = (nC_st1_b216_c0 == 0) ? nS_st1_b217_c0 : nS_st1_b217_c1;
  assign nS_st2_b218_c0 = nS_st1_b218_c0;
  assign nS_st2_b219_c0 = (nC_st1_b218_c0 == 0) ? nS_st1_b219_c0 : nS_st1_b219_c1;
  assign nS_st2_b220_c0 = nS_st1_b220_c0;
  assign nS_st2_b221_c0 = (nC_st1_b220_c0 == 0) ? nS_st1_b221_c0 : nS_st1_b221_c1;
  assign nS_st2_b222_c0 = nS_st1_b222_c0;
  assign nS_st2_b223_c0 = (nC_st1_b222_c0 == 0) ? nS_st1_b223_c0 : nS_st1_b223_c1;
  assign nS_st2_b224_c0 = nS_st1_b224_c0;
  assign nS_st2_b225_c0 = (nC_st1_b224_c0 == 0) ? nS_st1_b225_c0 : nS_st1_b225_c1;
  assign nS_st2_b226_c0 = nS_st1_b226_c0;
  assign nS_st2_b227_c0 = (nC_st1_b226_c0 == 0) ? nS_st1_b227_c0 : nS_st1_b227_c1;
  assign nS_st2_b228_c0 = nS_st1_b228_c0;
  assign nS_st2_b229_c0 = (nC_st1_b228_c0 == 0) ? nS_st1_b229_c0 : nS_st1_b229_c1;
  assign nS_st2_b230_c0 = nS_st1_b230_c0;
  assign nS_st2_b231_c0 = (nC_st1_b230_c0 == 0) ? nS_st1_b231_c0 : nS_st1_b231_c1;
  assign nS_st2_b232_c0 = nS_st1_b232_c0;
  assign nS_st2_b233_c0 = (nC_st1_b232_c0 == 0) ? nS_st1_b233_c0 : nS_st1_b233_c1;
  assign nS_st2_b234_c0 = nS_st1_b234_c0;
  assign nS_st2_b235_c0 = (nC_st1_b234_c0 == 0) ? nS_st1_b235_c0 : nS_st1_b235_c1;
  assign nS_st2_b236_c0 = nS_st1_b236_c0;
  assign nS_st2_b237_c0 = (nC_st1_b236_c0 == 0) ? nS_st1_b237_c0 : nS_st1_b237_c1;
  assign nS_st2_b238_c0 = nS_st1_b238_c0;
  assign nS_st2_b239_c0 = (nC_st1_b238_c0 == 0) ? nS_st1_b239_c0 : nS_st1_b239_c1;
  assign nS_st2_b240_c0 = nS_st1_b240_c0;
  assign nS_st2_b241_c0 = (nC_st1_b240_c0 == 0) ? nS_st1_b241_c0 : nS_st1_b241_c1;
  assign nS_st2_b242_c0 = nS_st1_b242_c0;
  assign nS_st2_b243_c0 = (nC_st1_b242_c0 == 0) ? nS_st1_b243_c0 : nS_st1_b243_c1;
  assign nS_st2_b244_c0 = nS_st1_b244_c0;
  assign nS_st2_b245_c0 = (nC_st1_b244_c0 == 0) ? nS_st1_b245_c0 : nS_st1_b245_c1;
  assign nS_st2_b246_c0 = nS_st1_b246_c0;
  assign nS_st2_b247_c0 = (nC_st1_b246_c0 == 0) ? nS_st1_b247_c0 : nS_st1_b247_c1;
  assign nS_st2_b248_c0 = nS_st1_b248_c0;
  assign nS_st2_b249_c0 = (nC_st1_b248_c0 == 0) ? nS_st1_b249_c0 : nS_st1_b249_c1;
  assign nS_st2_b250_c0 = nS_st1_b250_c0;
  assign nS_st2_b251_c0 = (nC_st1_b250_c0 == 0) ? nS_st1_b251_c0 : nS_st1_b251_c1;
  assign nS_st2_b252_c0 = nS_st1_b252_c0;
  assign nS_st2_b253_c0 = (nC_st1_b252_c0 == 0) ? nS_st1_b253_c0 : nS_st1_b253_c1;
  assign nS_st2_b254_c0 = nS_st1_b254_c0;
  assign nS_st2_b255_c0 = (nC_st1_b254_c0 == 0) ? nS_st1_b255_c0 : nS_st1_b255_c1;
  assign nS_st2_b0_c1 = nS_st1_b0_c1;
  assign nS_st2_b1_c1 = (nC_st1_b0_c1 == 0) ? nS_st1_b1_c0 : nS_st1_b1_c1;
  assign nS_st2_b2_c1 = nS_st1_b2_c1;
  assign nS_st2_b3_c1 = (nC_st1_b2_c1 == 0) ? nS_st1_b3_c0 : nS_st1_b3_c1;
  assign nS_st2_b4_c1 = nS_st1_b4_c1;
  assign nS_st2_b5_c1 = (nC_st1_b4_c1 == 0) ? nS_st1_b5_c0 : nS_st1_b5_c1;
  assign nS_st2_b6_c1 = nS_st1_b6_c1;
  assign nS_st2_b7_c1 = (nC_st1_b6_c1 == 0) ? nS_st1_b7_c0 : nS_st1_b7_c1;
  assign nS_st2_b8_c1 = nS_st1_b8_c1;
  assign nS_st2_b9_c1 = (nC_st1_b8_c1 == 0) ? nS_st1_b9_c0 : nS_st1_b9_c1;
  assign nS_st2_b10_c1 = nS_st1_b10_c1;
  assign nS_st2_b11_c1 = (nC_st1_b10_c1 == 0) ? nS_st1_b11_c0 : nS_st1_b11_c1;
  assign nS_st2_b12_c1 = nS_st1_b12_c1;
  assign nS_st2_b13_c1 = (nC_st1_b12_c1 == 0) ? nS_st1_b13_c0 : nS_st1_b13_c1;
  assign nS_st2_b14_c1 = nS_st1_b14_c1;
  assign nS_st2_b15_c1 = (nC_st1_b14_c1 == 0) ? nS_st1_b15_c0 : nS_st1_b15_c1;
  assign nS_st2_b16_c1 = nS_st1_b16_c1;
  assign nS_st2_b17_c1 = (nC_st1_b16_c1 == 0) ? nS_st1_b17_c0 : nS_st1_b17_c1;
  assign nS_st2_b18_c1 = nS_st1_b18_c1;
  assign nS_st2_b19_c1 = (nC_st1_b18_c1 == 0) ? nS_st1_b19_c0 : nS_st1_b19_c1;
  assign nS_st2_b20_c1 = nS_st1_b20_c1;
  assign nS_st2_b21_c1 = (nC_st1_b20_c1 == 0) ? nS_st1_b21_c0 : nS_st1_b21_c1;
  assign nS_st2_b22_c1 = nS_st1_b22_c1;
  assign nS_st2_b23_c1 = (nC_st1_b22_c1 == 0) ? nS_st1_b23_c0 : nS_st1_b23_c1;
  assign nS_st2_b24_c1 = nS_st1_b24_c1;
  assign nS_st2_b25_c1 = (nC_st1_b24_c1 == 0) ? nS_st1_b25_c0 : nS_st1_b25_c1;
  assign nS_st2_b26_c1 = nS_st1_b26_c1;
  assign nS_st2_b27_c1 = (nC_st1_b26_c1 == 0) ? nS_st1_b27_c0 : nS_st1_b27_c1;
  assign nS_st2_b28_c1 = nS_st1_b28_c1;
  assign nS_st2_b29_c1 = (nC_st1_b28_c1 == 0) ? nS_st1_b29_c0 : nS_st1_b29_c1;
  assign nS_st2_b30_c1 = nS_st1_b30_c1;
  assign nS_st2_b31_c1 = (nC_st1_b30_c1 == 0) ? nS_st1_b31_c0 : nS_st1_b31_c1;
  assign nS_st2_b32_c1 = nS_st1_b32_c1;
  assign nS_st2_b33_c1 = (nC_st1_b32_c1 == 0) ? nS_st1_b33_c0 : nS_st1_b33_c1;
  assign nS_st2_b34_c1 = nS_st1_b34_c1;
  assign nS_st2_b35_c1 = (nC_st1_b34_c1 == 0) ? nS_st1_b35_c0 : nS_st1_b35_c1;
  assign nS_st2_b36_c1 = nS_st1_b36_c1;
  assign nS_st2_b37_c1 = (nC_st1_b36_c1 == 0) ? nS_st1_b37_c0 : nS_st1_b37_c1;
  assign nS_st2_b38_c1 = nS_st1_b38_c1;
  assign nS_st2_b39_c1 = (nC_st1_b38_c1 == 0) ? nS_st1_b39_c0 : nS_st1_b39_c1;
  assign nS_st2_b40_c1 = nS_st1_b40_c1;
  assign nS_st2_b41_c1 = (nC_st1_b40_c1 == 0) ? nS_st1_b41_c0 : nS_st1_b41_c1;
  assign nS_st2_b42_c1 = nS_st1_b42_c1;
  assign nS_st2_b43_c1 = (nC_st1_b42_c1 == 0) ? nS_st1_b43_c0 : nS_st1_b43_c1;
  assign nS_st2_b44_c1 = nS_st1_b44_c1;
  assign nS_st2_b45_c1 = (nC_st1_b44_c1 == 0) ? nS_st1_b45_c0 : nS_st1_b45_c1;
  assign nS_st2_b46_c1 = nS_st1_b46_c1;
  assign nS_st2_b47_c1 = (nC_st1_b46_c1 == 0) ? nS_st1_b47_c0 : nS_st1_b47_c1;
  assign nS_st2_b48_c1 = nS_st1_b48_c1;
  assign nS_st2_b49_c1 = (nC_st1_b48_c1 == 0) ? nS_st1_b49_c0 : nS_st1_b49_c1;
  assign nS_st2_b50_c1 = nS_st1_b50_c1;
  assign nS_st2_b51_c1 = (nC_st1_b50_c1 == 0) ? nS_st1_b51_c0 : nS_st1_b51_c1;
  assign nS_st2_b52_c1 = nS_st1_b52_c1;
  assign nS_st2_b53_c1 = (nC_st1_b52_c1 == 0) ? nS_st1_b53_c0 : nS_st1_b53_c1;
  assign nS_st2_b54_c1 = nS_st1_b54_c1;
  assign nS_st2_b55_c1 = (nC_st1_b54_c1 == 0) ? nS_st1_b55_c0 : nS_st1_b55_c1;
  assign nS_st2_b56_c1 = nS_st1_b56_c1;
  assign nS_st2_b57_c1 = (nC_st1_b56_c1 == 0) ? nS_st1_b57_c0 : nS_st1_b57_c1;
  assign nS_st2_b58_c1 = nS_st1_b58_c1;
  assign nS_st2_b59_c1 = (nC_st1_b58_c1 == 0) ? nS_st1_b59_c0 : nS_st1_b59_c1;
  assign nS_st2_b60_c1 = nS_st1_b60_c1;
  assign nS_st2_b61_c1 = (nC_st1_b60_c1 == 0) ? nS_st1_b61_c0 : nS_st1_b61_c1;
  assign nS_st2_b62_c1 = nS_st1_b62_c1;
  assign nS_st2_b63_c1 = (nC_st1_b62_c1 == 0) ? nS_st1_b63_c0 : nS_st1_b63_c1;
  assign nS_st2_b64_c1 = nS_st1_b64_c1;
  assign nS_st2_b65_c1 = (nC_st1_b64_c1 == 0) ? nS_st1_b65_c0 : nS_st1_b65_c1;
  assign nS_st2_b66_c1 = nS_st1_b66_c1;
  assign nS_st2_b67_c1 = (nC_st1_b66_c1 == 0) ? nS_st1_b67_c0 : nS_st1_b67_c1;
  assign nS_st2_b68_c1 = nS_st1_b68_c1;
  assign nS_st2_b69_c1 = (nC_st1_b68_c1 == 0) ? nS_st1_b69_c0 : nS_st1_b69_c1;
  assign nS_st2_b70_c1 = nS_st1_b70_c1;
  assign nS_st2_b71_c1 = (nC_st1_b70_c1 == 0) ? nS_st1_b71_c0 : nS_st1_b71_c1;
  assign nS_st2_b72_c1 = nS_st1_b72_c1;
  assign nS_st2_b73_c1 = (nC_st1_b72_c1 == 0) ? nS_st1_b73_c0 : nS_st1_b73_c1;
  assign nS_st2_b74_c1 = nS_st1_b74_c1;
  assign nS_st2_b75_c1 = (nC_st1_b74_c1 == 0) ? nS_st1_b75_c0 : nS_st1_b75_c1;
  assign nS_st2_b76_c1 = nS_st1_b76_c1;
  assign nS_st2_b77_c1 = (nC_st1_b76_c1 == 0) ? nS_st1_b77_c0 : nS_st1_b77_c1;
  assign nS_st2_b78_c1 = nS_st1_b78_c1;
  assign nS_st2_b79_c1 = (nC_st1_b78_c1 == 0) ? nS_st1_b79_c0 : nS_st1_b79_c1;
  assign nS_st2_b80_c1 = nS_st1_b80_c1;
  assign nS_st2_b81_c1 = (nC_st1_b80_c1 == 0) ? nS_st1_b81_c0 : nS_st1_b81_c1;
  assign nS_st2_b82_c1 = nS_st1_b82_c1;
  assign nS_st2_b83_c1 = (nC_st1_b82_c1 == 0) ? nS_st1_b83_c0 : nS_st1_b83_c1;
  assign nS_st2_b84_c1 = nS_st1_b84_c1;
  assign nS_st2_b85_c1 = (nC_st1_b84_c1 == 0) ? nS_st1_b85_c0 : nS_st1_b85_c1;
  assign nS_st2_b86_c1 = nS_st1_b86_c1;
  assign nS_st2_b87_c1 = (nC_st1_b86_c1 == 0) ? nS_st1_b87_c0 : nS_st1_b87_c1;
  assign nS_st2_b88_c1 = nS_st1_b88_c1;
  assign nS_st2_b89_c1 = (nC_st1_b88_c1 == 0) ? nS_st1_b89_c0 : nS_st1_b89_c1;
  assign nS_st2_b90_c1 = nS_st1_b90_c1;
  assign nS_st2_b91_c1 = (nC_st1_b90_c1 == 0) ? nS_st1_b91_c0 : nS_st1_b91_c1;
  assign nS_st2_b92_c1 = nS_st1_b92_c1;
  assign nS_st2_b93_c1 = (nC_st1_b92_c1 == 0) ? nS_st1_b93_c0 : nS_st1_b93_c1;
  assign nS_st2_b94_c1 = nS_st1_b94_c1;
  assign nS_st2_b95_c1 = (nC_st1_b94_c1 == 0) ? nS_st1_b95_c0 : nS_st1_b95_c1;
  assign nS_st2_b96_c1 = nS_st1_b96_c1;
  assign nS_st2_b97_c1 = (nC_st1_b96_c1 == 0) ? nS_st1_b97_c0 : nS_st1_b97_c1;
  assign nS_st2_b98_c1 = nS_st1_b98_c1;
  assign nS_st2_b99_c1 = (nC_st1_b98_c1 == 0) ? nS_st1_b99_c0 : nS_st1_b99_c1;
  assign nS_st2_b100_c1 = nS_st1_b100_c1;
  assign nS_st2_b101_c1 = (nC_st1_b100_c1 == 0) ? nS_st1_b101_c0 : nS_st1_b101_c1;
  assign nS_st2_b102_c1 = nS_st1_b102_c1;
  assign nS_st2_b103_c1 = (nC_st1_b102_c1 == 0) ? nS_st1_b103_c0 : nS_st1_b103_c1;
  assign nS_st2_b104_c1 = nS_st1_b104_c1;
  assign nS_st2_b105_c1 = (nC_st1_b104_c1 == 0) ? nS_st1_b105_c0 : nS_st1_b105_c1;
  assign nS_st2_b106_c1 = nS_st1_b106_c1;
  assign nS_st2_b107_c1 = (nC_st1_b106_c1 == 0) ? nS_st1_b107_c0 : nS_st1_b107_c1;
  assign nS_st2_b108_c1 = nS_st1_b108_c1;
  assign nS_st2_b109_c1 = (nC_st1_b108_c1 == 0) ? nS_st1_b109_c0 : nS_st1_b109_c1;
  assign nS_st2_b110_c1 = nS_st1_b110_c1;
  assign nS_st2_b111_c1 = (nC_st1_b110_c1 == 0) ? nS_st1_b111_c0 : nS_st1_b111_c1;
  assign nS_st2_b112_c1 = nS_st1_b112_c1;
  assign nS_st2_b113_c1 = (nC_st1_b112_c1 == 0) ? nS_st1_b113_c0 : nS_st1_b113_c1;
  assign nS_st2_b114_c1 = nS_st1_b114_c1;
  assign nS_st2_b115_c1 = (nC_st1_b114_c1 == 0) ? nS_st1_b115_c0 : nS_st1_b115_c1;
  assign nS_st2_b116_c1 = nS_st1_b116_c1;
  assign nS_st2_b117_c1 = (nC_st1_b116_c1 == 0) ? nS_st1_b117_c0 : nS_st1_b117_c1;
  assign nS_st2_b118_c1 = nS_st1_b118_c1;
  assign nS_st2_b119_c1 = (nC_st1_b118_c1 == 0) ? nS_st1_b119_c0 : nS_st1_b119_c1;
  assign nS_st2_b120_c1 = nS_st1_b120_c1;
  assign nS_st2_b121_c1 = (nC_st1_b120_c1 == 0) ? nS_st1_b121_c0 : nS_st1_b121_c1;
  assign nS_st2_b122_c1 = nS_st1_b122_c1;
  assign nS_st2_b123_c1 = (nC_st1_b122_c1 == 0) ? nS_st1_b123_c0 : nS_st1_b123_c1;
  assign nS_st2_b124_c1 = nS_st1_b124_c1;
  assign nS_st2_b125_c1 = (nC_st1_b124_c1 == 0) ? nS_st1_b125_c0 : nS_st1_b125_c1;
  assign nS_st2_b126_c1 = nS_st1_b126_c1;
  assign nS_st2_b127_c1 = (nC_st1_b126_c1 == 0) ? nS_st1_b127_c0 : nS_st1_b127_c1;
  assign nS_st2_b128_c1 = nS_st1_b128_c1;
  assign nS_st2_b129_c1 = (nC_st1_b128_c1 == 0) ? nS_st1_b129_c0 : nS_st1_b129_c1;
  assign nS_st2_b130_c1 = nS_st1_b130_c1;
  assign nS_st2_b131_c1 = (nC_st1_b130_c1 == 0) ? nS_st1_b131_c0 : nS_st1_b131_c1;
  assign nS_st2_b132_c1 = nS_st1_b132_c1;
  assign nS_st2_b133_c1 = (nC_st1_b132_c1 == 0) ? nS_st1_b133_c0 : nS_st1_b133_c1;
  assign nS_st2_b134_c1 = nS_st1_b134_c1;
  assign nS_st2_b135_c1 = (nC_st1_b134_c1 == 0) ? nS_st1_b135_c0 : nS_st1_b135_c1;
  assign nS_st2_b136_c1 = nS_st1_b136_c1;
  assign nS_st2_b137_c1 = (nC_st1_b136_c1 == 0) ? nS_st1_b137_c0 : nS_st1_b137_c1;
  assign nS_st2_b138_c1 = nS_st1_b138_c1;
  assign nS_st2_b139_c1 = (nC_st1_b138_c1 == 0) ? nS_st1_b139_c0 : nS_st1_b139_c1;
  assign nS_st2_b140_c1 = nS_st1_b140_c1;
  assign nS_st2_b141_c1 = (nC_st1_b140_c1 == 0) ? nS_st1_b141_c0 : nS_st1_b141_c1;
  assign nS_st2_b142_c1 = nS_st1_b142_c1;
  assign nS_st2_b143_c1 = (nC_st1_b142_c1 == 0) ? nS_st1_b143_c0 : nS_st1_b143_c1;
  assign nS_st2_b144_c1 = nS_st1_b144_c1;
  assign nS_st2_b145_c1 = (nC_st1_b144_c1 == 0) ? nS_st1_b145_c0 : nS_st1_b145_c1;
  assign nS_st2_b146_c1 = nS_st1_b146_c1;
  assign nS_st2_b147_c1 = (nC_st1_b146_c1 == 0) ? nS_st1_b147_c0 : nS_st1_b147_c1;
  assign nS_st2_b148_c1 = nS_st1_b148_c1;
  assign nS_st2_b149_c1 = (nC_st1_b148_c1 == 0) ? nS_st1_b149_c0 : nS_st1_b149_c1;
  assign nS_st2_b150_c1 = nS_st1_b150_c1;
  assign nS_st2_b151_c1 = (nC_st1_b150_c1 == 0) ? nS_st1_b151_c0 : nS_st1_b151_c1;
  assign nS_st2_b152_c1 = nS_st1_b152_c1;
  assign nS_st2_b153_c1 = (nC_st1_b152_c1 == 0) ? nS_st1_b153_c0 : nS_st1_b153_c1;
  assign nS_st2_b154_c1 = nS_st1_b154_c1;
  assign nS_st2_b155_c1 = (nC_st1_b154_c1 == 0) ? nS_st1_b155_c0 : nS_st1_b155_c1;
  assign nS_st2_b156_c1 = nS_st1_b156_c1;
  assign nS_st2_b157_c1 = (nC_st1_b156_c1 == 0) ? nS_st1_b157_c0 : nS_st1_b157_c1;
  assign nS_st2_b158_c1 = nS_st1_b158_c1;
  assign nS_st2_b159_c1 = (nC_st1_b158_c1 == 0) ? nS_st1_b159_c0 : nS_st1_b159_c1;
  assign nS_st2_b160_c1 = nS_st1_b160_c1;
  assign nS_st2_b161_c1 = (nC_st1_b160_c1 == 0) ? nS_st1_b161_c0 : nS_st1_b161_c1;
  assign nS_st2_b162_c1 = nS_st1_b162_c1;
  assign nS_st2_b163_c1 = (nC_st1_b162_c1 == 0) ? nS_st1_b163_c0 : nS_st1_b163_c1;
  assign nS_st2_b164_c1 = nS_st1_b164_c1;
  assign nS_st2_b165_c1 = (nC_st1_b164_c1 == 0) ? nS_st1_b165_c0 : nS_st1_b165_c1;
  assign nS_st2_b166_c1 = nS_st1_b166_c1;
  assign nS_st2_b167_c1 = (nC_st1_b166_c1 == 0) ? nS_st1_b167_c0 : nS_st1_b167_c1;
  assign nS_st2_b168_c1 = nS_st1_b168_c1;
  assign nS_st2_b169_c1 = (nC_st1_b168_c1 == 0) ? nS_st1_b169_c0 : nS_st1_b169_c1;
  assign nS_st2_b170_c1 = nS_st1_b170_c1;
  assign nS_st2_b171_c1 = (nC_st1_b170_c1 == 0) ? nS_st1_b171_c0 : nS_st1_b171_c1;
  assign nS_st2_b172_c1 = nS_st1_b172_c1;
  assign nS_st2_b173_c1 = (nC_st1_b172_c1 == 0) ? nS_st1_b173_c0 : nS_st1_b173_c1;
  assign nS_st2_b174_c1 = nS_st1_b174_c1;
  assign nS_st2_b175_c1 = (nC_st1_b174_c1 == 0) ? nS_st1_b175_c0 : nS_st1_b175_c1;
  assign nS_st2_b176_c1 = nS_st1_b176_c1;
  assign nS_st2_b177_c1 = (nC_st1_b176_c1 == 0) ? nS_st1_b177_c0 : nS_st1_b177_c1;
  assign nS_st2_b178_c1 = nS_st1_b178_c1;
  assign nS_st2_b179_c1 = (nC_st1_b178_c1 == 0) ? nS_st1_b179_c0 : nS_st1_b179_c1;
  assign nS_st2_b180_c1 = nS_st1_b180_c1;
  assign nS_st2_b181_c1 = (nC_st1_b180_c1 == 0) ? nS_st1_b181_c0 : nS_st1_b181_c1;
  assign nS_st2_b182_c1 = nS_st1_b182_c1;
  assign nS_st2_b183_c1 = (nC_st1_b182_c1 == 0) ? nS_st1_b183_c0 : nS_st1_b183_c1;
  assign nS_st2_b184_c1 = nS_st1_b184_c1;
  assign nS_st2_b185_c1 = (nC_st1_b184_c1 == 0) ? nS_st1_b185_c0 : nS_st1_b185_c1;
  assign nS_st2_b186_c1 = nS_st1_b186_c1;
  assign nS_st2_b187_c1 = (nC_st1_b186_c1 == 0) ? nS_st1_b187_c0 : nS_st1_b187_c1;
  assign nS_st2_b188_c1 = nS_st1_b188_c1;
  assign nS_st2_b189_c1 = (nC_st1_b188_c1 == 0) ? nS_st1_b189_c0 : nS_st1_b189_c1;
  assign nS_st2_b190_c1 = nS_st1_b190_c1;
  assign nS_st2_b191_c1 = (nC_st1_b190_c1 == 0) ? nS_st1_b191_c0 : nS_st1_b191_c1;
  assign nS_st2_b192_c1 = nS_st1_b192_c1;
  assign nS_st2_b193_c1 = (nC_st1_b192_c1 == 0) ? nS_st1_b193_c0 : nS_st1_b193_c1;
  assign nS_st2_b194_c1 = nS_st1_b194_c1;
  assign nS_st2_b195_c1 = (nC_st1_b194_c1 == 0) ? nS_st1_b195_c0 : nS_st1_b195_c1;
  assign nS_st2_b196_c1 = nS_st1_b196_c1;
  assign nS_st2_b197_c1 = (nC_st1_b196_c1 == 0) ? nS_st1_b197_c0 : nS_st1_b197_c1;
  assign nS_st2_b198_c1 = nS_st1_b198_c1;
  assign nS_st2_b199_c1 = (nC_st1_b198_c1 == 0) ? nS_st1_b199_c0 : nS_st1_b199_c1;
  assign nS_st2_b200_c1 = nS_st1_b200_c1;
  assign nS_st2_b201_c1 = (nC_st1_b200_c1 == 0) ? nS_st1_b201_c0 : nS_st1_b201_c1;
  assign nS_st2_b202_c1 = nS_st1_b202_c1;
  assign nS_st2_b203_c1 = (nC_st1_b202_c1 == 0) ? nS_st1_b203_c0 : nS_st1_b203_c1;
  assign nS_st2_b204_c1 = nS_st1_b204_c1;
  assign nS_st2_b205_c1 = (nC_st1_b204_c1 == 0) ? nS_st1_b205_c0 : nS_st1_b205_c1;
  assign nS_st2_b206_c1 = nS_st1_b206_c1;
  assign nS_st2_b207_c1 = (nC_st1_b206_c1 == 0) ? nS_st1_b207_c0 : nS_st1_b207_c1;
  assign nS_st2_b208_c1 = nS_st1_b208_c1;
  assign nS_st2_b209_c1 = (nC_st1_b208_c1 == 0) ? nS_st1_b209_c0 : nS_st1_b209_c1;
  assign nS_st2_b210_c1 = nS_st1_b210_c1;
  assign nS_st2_b211_c1 = (nC_st1_b210_c1 == 0) ? nS_st1_b211_c0 : nS_st1_b211_c1;
  assign nS_st2_b212_c1 = nS_st1_b212_c1;
  assign nS_st2_b213_c1 = (nC_st1_b212_c1 == 0) ? nS_st1_b213_c0 : nS_st1_b213_c1;
  assign nS_st2_b214_c1 = nS_st1_b214_c1;
  assign nS_st2_b215_c1 = (nC_st1_b214_c1 == 0) ? nS_st1_b215_c0 : nS_st1_b215_c1;
  assign nS_st2_b216_c1 = nS_st1_b216_c1;
  assign nS_st2_b217_c1 = (nC_st1_b216_c1 == 0) ? nS_st1_b217_c0 : nS_st1_b217_c1;
  assign nS_st2_b218_c1 = nS_st1_b218_c1;
  assign nS_st2_b219_c1 = (nC_st1_b218_c1 == 0) ? nS_st1_b219_c0 : nS_st1_b219_c1;
  assign nS_st2_b220_c1 = nS_st1_b220_c1;
  assign nS_st2_b221_c1 = (nC_st1_b220_c1 == 0) ? nS_st1_b221_c0 : nS_st1_b221_c1;
  assign nS_st2_b222_c1 = nS_st1_b222_c1;
  assign nS_st2_b223_c1 = (nC_st1_b222_c1 == 0) ? nS_st1_b223_c0 : nS_st1_b223_c1;
  assign nS_st2_b224_c1 = nS_st1_b224_c1;
  assign nS_st2_b225_c1 = (nC_st1_b224_c1 == 0) ? nS_st1_b225_c0 : nS_st1_b225_c1;
  assign nS_st2_b226_c1 = nS_st1_b226_c1;
  assign nS_st2_b227_c1 = (nC_st1_b226_c1 == 0) ? nS_st1_b227_c0 : nS_st1_b227_c1;
  assign nS_st2_b228_c1 = nS_st1_b228_c1;
  assign nS_st2_b229_c1 = (nC_st1_b228_c1 == 0) ? nS_st1_b229_c0 : nS_st1_b229_c1;
  assign nS_st2_b230_c1 = nS_st1_b230_c1;
  assign nS_st2_b231_c1 = (nC_st1_b230_c1 == 0) ? nS_st1_b231_c0 : nS_st1_b231_c1;
  assign nS_st2_b232_c1 = nS_st1_b232_c1;
  assign nS_st2_b233_c1 = (nC_st1_b232_c1 == 0) ? nS_st1_b233_c0 : nS_st1_b233_c1;
  assign nS_st2_b234_c1 = nS_st1_b234_c1;
  assign nS_st2_b235_c1 = (nC_st1_b234_c1 == 0) ? nS_st1_b235_c0 : nS_st1_b235_c1;
  assign nS_st2_b236_c1 = nS_st1_b236_c1;
  assign nS_st2_b237_c1 = (nC_st1_b236_c1 == 0) ? nS_st1_b237_c0 : nS_st1_b237_c1;
  assign nS_st2_b238_c1 = nS_st1_b238_c1;
  assign nS_st2_b239_c1 = (nC_st1_b238_c1 == 0) ? nS_st1_b239_c0 : nS_st1_b239_c1;
  assign nS_st2_b240_c1 = nS_st1_b240_c1;
  assign nS_st2_b241_c1 = (nC_st1_b240_c1 == 0) ? nS_st1_b241_c0 : nS_st1_b241_c1;
  assign nS_st2_b242_c1 = nS_st1_b242_c1;
  assign nS_st2_b243_c1 = (nC_st1_b242_c1 == 0) ? nS_st1_b243_c0 : nS_st1_b243_c1;
  assign nS_st2_b244_c1 = nS_st1_b244_c1;
  assign nS_st2_b245_c1 = (nC_st1_b244_c1 == 0) ? nS_st1_b245_c0 : nS_st1_b245_c1;
  assign nS_st2_b246_c1 = nS_st1_b246_c1;
  assign nS_st2_b247_c1 = (nC_st1_b246_c1 == 0) ? nS_st1_b247_c0 : nS_st1_b247_c1;
  assign nS_st2_b248_c1 = nS_st1_b248_c1;
  assign nS_st2_b249_c1 = (nC_st1_b248_c1 == 0) ? nS_st1_b249_c0 : nS_st1_b249_c1;
  assign nS_st2_b250_c1 = nS_st1_b250_c1;
  assign nS_st2_b251_c1 = (nC_st1_b250_c1 == 0) ? nS_st1_b251_c0 : nS_st1_b251_c1;
  assign nS_st2_b252_c1 = nS_st1_b252_c1;
  assign nS_st2_b253_c1 = (nC_st1_b252_c1 == 0) ? nS_st1_b253_c0 : nS_st1_b253_c1;
  assign nS_st2_b254_c1 = nS_st1_b254_c1;
  assign nS_st2_b255_c1 = (nC_st1_b254_c1 == 0) ? nS_st1_b255_c0 : nS_st1_b255_c1;
  assign nC_st2_b1_c0 = (nC_st1_b0_c0 == 0) ? nC_st1_b1_c0 : nC_st1_b1_c1;
  assign nC_st2_b3_c0 = (nC_st1_b2_c0 == 0) ? nC_st1_b3_c0 : nC_st1_b3_c1;
  assign nC_st2_b5_c0 = (nC_st1_b4_c0 == 0) ? nC_st1_b5_c0 : nC_st1_b5_c1;
  assign nC_st2_b7_c0 = (nC_st1_b6_c0 == 0) ? nC_st1_b7_c0 : nC_st1_b7_c1;
  assign nC_st2_b9_c0 = (nC_st1_b8_c0 == 0) ? nC_st1_b9_c0 : nC_st1_b9_c1;
  assign nC_st2_b11_c0 = (nC_st1_b10_c0 == 0) ? nC_st1_b11_c0 : nC_st1_b11_c1;
  assign nC_st2_b13_c0 = (nC_st1_b12_c0 == 0) ? nC_st1_b13_c0 : nC_st1_b13_c1;
  assign nC_st2_b15_c0 = (nC_st1_b14_c0 == 0) ? nC_st1_b15_c0 : nC_st1_b15_c1;
  assign nC_st2_b17_c0 = (nC_st1_b16_c0 == 0) ? nC_st1_b17_c0 : nC_st1_b17_c1;
  assign nC_st2_b19_c0 = (nC_st1_b18_c0 == 0) ? nC_st1_b19_c0 : nC_st1_b19_c1;
  assign nC_st2_b21_c0 = (nC_st1_b20_c0 == 0) ? nC_st1_b21_c0 : nC_st1_b21_c1;
  assign nC_st2_b23_c0 = (nC_st1_b22_c0 == 0) ? nC_st1_b23_c0 : nC_st1_b23_c1;
  assign nC_st2_b25_c0 = (nC_st1_b24_c0 == 0) ? nC_st1_b25_c0 : nC_st1_b25_c1;
  assign nC_st2_b27_c0 = (nC_st1_b26_c0 == 0) ? nC_st1_b27_c0 : nC_st1_b27_c1;
  assign nC_st2_b29_c0 = (nC_st1_b28_c0 == 0) ? nC_st1_b29_c0 : nC_st1_b29_c1;
  assign nC_st2_b31_c0 = (nC_st1_b30_c0 == 0) ? nC_st1_b31_c0 : nC_st1_b31_c1;
  assign nC_st2_b33_c0 = (nC_st1_b32_c0 == 0) ? nC_st1_b33_c0 : nC_st1_b33_c1;
  assign nC_st2_b35_c0 = (nC_st1_b34_c0 == 0) ? nC_st1_b35_c0 : nC_st1_b35_c1;
  assign nC_st2_b37_c0 = (nC_st1_b36_c0 == 0) ? nC_st1_b37_c0 : nC_st1_b37_c1;
  assign nC_st2_b39_c0 = (nC_st1_b38_c0 == 0) ? nC_st1_b39_c0 : nC_st1_b39_c1;
  assign nC_st2_b41_c0 = (nC_st1_b40_c0 == 0) ? nC_st1_b41_c0 : nC_st1_b41_c1;
  assign nC_st2_b43_c0 = (nC_st1_b42_c0 == 0) ? nC_st1_b43_c0 : nC_st1_b43_c1;
  assign nC_st2_b45_c0 = (nC_st1_b44_c0 == 0) ? nC_st1_b45_c0 : nC_st1_b45_c1;
  assign nC_st2_b47_c0 = (nC_st1_b46_c0 == 0) ? nC_st1_b47_c0 : nC_st1_b47_c1;
  assign nC_st2_b49_c0 = (nC_st1_b48_c0 == 0) ? nC_st1_b49_c0 : nC_st1_b49_c1;
  assign nC_st2_b51_c0 = (nC_st1_b50_c0 == 0) ? nC_st1_b51_c0 : nC_st1_b51_c1;
  assign nC_st2_b53_c0 = (nC_st1_b52_c0 == 0) ? nC_st1_b53_c0 : nC_st1_b53_c1;
  assign nC_st2_b55_c0 = (nC_st1_b54_c0 == 0) ? nC_st1_b55_c0 : nC_st1_b55_c1;
  assign nC_st2_b57_c0 = (nC_st1_b56_c0 == 0) ? nC_st1_b57_c0 : nC_st1_b57_c1;
  assign nC_st2_b59_c0 = (nC_st1_b58_c0 == 0) ? nC_st1_b59_c0 : nC_st1_b59_c1;
  assign nC_st2_b61_c0 = (nC_st1_b60_c0 == 0) ? nC_st1_b61_c0 : nC_st1_b61_c1;
  assign nC_st2_b63_c0 = (nC_st1_b62_c0 == 0) ? nC_st1_b63_c0 : nC_st1_b63_c1;
  assign nC_st2_b65_c0 = (nC_st1_b64_c0 == 0) ? nC_st1_b65_c0 : nC_st1_b65_c1;
  assign nC_st2_b67_c0 = (nC_st1_b66_c0 == 0) ? nC_st1_b67_c0 : nC_st1_b67_c1;
  assign nC_st2_b69_c0 = (nC_st1_b68_c0 == 0) ? nC_st1_b69_c0 : nC_st1_b69_c1;
  assign nC_st2_b71_c0 = (nC_st1_b70_c0 == 0) ? nC_st1_b71_c0 : nC_st1_b71_c1;
  assign nC_st2_b73_c0 = (nC_st1_b72_c0 == 0) ? nC_st1_b73_c0 : nC_st1_b73_c1;
  assign nC_st2_b75_c0 = (nC_st1_b74_c0 == 0) ? nC_st1_b75_c0 : nC_st1_b75_c1;
  assign nC_st2_b77_c0 = (nC_st1_b76_c0 == 0) ? nC_st1_b77_c0 : nC_st1_b77_c1;
  assign nC_st2_b79_c0 = (nC_st1_b78_c0 == 0) ? nC_st1_b79_c0 : nC_st1_b79_c1;
  assign nC_st2_b81_c0 = (nC_st1_b80_c0 == 0) ? nC_st1_b81_c0 : nC_st1_b81_c1;
  assign nC_st2_b83_c0 = (nC_st1_b82_c0 == 0) ? nC_st1_b83_c0 : nC_st1_b83_c1;
  assign nC_st2_b85_c0 = (nC_st1_b84_c0 == 0) ? nC_st1_b85_c0 : nC_st1_b85_c1;
  assign nC_st2_b87_c0 = (nC_st1_b86_c0 == 0) ? nC_st1_b87_c0 : nC_st1_b87_c1;
  assign nC_st2_b89_c0 = (nC_st1_b88_c0 == 0) ? nC_st1_b89_c0 : nC_st1_b89_c1;
  assign nC_st2_b91_c0 = (nC_st1_b90_c0 == 0) ? nC_st1_b91_c0 : nC_st1_b91_c1;
  assign nC_st2_b93_c0 = (nC_st1_b92_c0 == 0) ? nC_st1_b93_c0 : nC_st1_b93_c1;
  assign nC_st2_b95_c0 = (nC_st1_b94_c0 == 0) ? nC_st1_b95_c0 : nC_st1_b95_c1;
  assign nC_st2_b97_c0 = (nC_st1_b96_c0 == 0) ? nC_st1_b97_c0 : nC_st1_b97_c1;
  assign nC_st2_b99_c0 = (nC_st1_b98_c0 == 0) ? nC_st1_b99_c0 : nC_st1_b99_c1;
  assign nC_st2_b101_c0 = (nC_st1_b100_c0 == 0) ? nC_st1_b101_c0 : nC_st1_b101_c1;
  assign nC_st2_b103_c0 = (nC_st1_b102_c0 == 0) ? nC_st1_b103_c0 : nC_st1_b103_c1;
  assign nC_st2_b105_c0 = (nC_st1_b104_c0 == 0) ? nC_st1_b105_c0 : nC_st1_b105_c1;
  assign nC_st2_b107_c0 = (nC_st1_b106_c0 == 0) ? nC_st1_b107_c0 : nC_st1_b107_c1;
  assign nC_st2_b109_c0 = (nC_st1_b108_c0 == 0) ? nC_st1_b109_c0 : nC_st1_b109_c1;
  assign nC_st2_b111_c0 = (nC_st1_b110_c0 == 0) ? nC_st1_b111_c0 : nC_st1_b111_c1;
  assign nC_st2_b113_c0 = (nC_st1_b112_c0 == 0) ? nC_st1_b113_c0 : nC_st1_b113_c1;
  assign nC_st2_b115_c0 = (nC_st1_b114_c0 == 0) ? nC_st1_b115_c0 : nC_st1_b115_c1;
  assign nC_st2_b117_c0 = (nC_st1_b116_c0 == 0) ? nC_st1_b117_c0 : nC_st1_b117_c1;
  assign nC_st2_b119_c0 = (nC_st1_b118_c0 == 0) ? nC_st1_b119_c0 : nC_st1_b119_c1;
  assign nC_st2_b121_c0 = (nC_st1_b120_c0 == 0) ? nC_st1_b121_c0 : nC_st1_b121_c1;
  assign nC_st2_b123_c0 = (nC_st1_b122_c0 == 0) ? nC_st1_b123_c0 : nC_st1_b123_c1;
  assign nC_st2_b125_c0 = (nC_st1_b124_c0 == 0) ? nC_st1_b125_c0 : nC_st1_b125_c1;
  assign nC_st2_b127_c0 = (nC_st1_b126_c0 == 0) ? nC_st1_b127_c0 : nC_st1_b127_c1;
  assign nC_st2_b129_c0 = (nC_st1_b128_c0 == 0) ? nC_st1_b129_c0 : nC_st1_b129_c1;
  assign nC_st2_b131_c0 = (nC_st1_b130_c0 == 0) ? nC_st1_b131_c0 : nC_st1_b131_c1;
  assign nC_st2_b133_c0 = (nC_st1_b132_c0 == 0) ? nC_st1_b133_c0 : nC_st1_b133_c1;
  assign nC_st2_b135_c0 = (nC_st1_b134_c0 == 0) ? nC_st1_b135_c0 : nC_st1_b135_c1;
  assign nC_st2_b137_c0 = (nC_st1_b136_c0 == 0) ? nC_st1_b137_c0 : nC_st1_b137_c1;
  assign nC_st2_b139_c0 = (nC_st1_b138_c0 == 0) ? nC_st1_b139_c0 : nC_st1_b139_c1;
  assign nC_st2_b141_c0 = (nC_st1_b140_c0 == 0) ? nC_st1_b141_c0 : nC_st1_b141_c1;
  assign nC_st2_b143_c0 = (nC_st1_b142_c0 == 0) ? nC_st1_b143_c0 : nC_st1_b143_c1;
  assign nC_st2_b145_c0 = (nC_st1_b144_c0 == 0) ? nC_st1_b145_c0 : nC_st1_b145_c1;
  assign nC_st2_b147_c0 = (nC_st1_b146_c0 == 0) ? nC_st1_b147_c0 : nC_st1_b147_c1;
  assign nC_st2_b149_c0 = (nC_st1_b148_c0 == 0) ? nC_st1_b149_c0 : nC_st1_b149_c1;
  assign nC_st2_b151_c0 = (nC_st1_b150_c0 == 0) ? nC_st1_b151_c0 : nC_st1_b151_c1;
  assign nC_st2_b153_c0 = (nC_st1_b152_c0 == 0) ? nC_st1_b153_c0 : nC_st1_b153_c1;
  assign nC_st2_b155_c0 = (nC_st1_b154_c0 == 0) ? nC_st1_b155_c0 : nC_st1_b155_c1;
  assign nC_st2_b157_c0 = (nC_st1_b156_c0 == 0) ? nC_st1_b157_c0 : nC_st1_b157_c1;
  assign nC_st2_b159_c0 = (nC_st1_b158_c0 == 0) ? nC_st1_b159_c0 : nC_st1_b159_c1;
  assign nC_st2_b161_c0 = (nC_st1_b160_c0 == 0) ? nC_st1_b161_c0 : nC_st1_b161_c1;
  assign nC_st2_b163_c0 = (nC_st1_b162_c0 == 0) ? nC_st1_b163_c0 : nC_st1_b163_c1;
  assign nC_st2_b165_c0 = (nC_st1_b164_c0 == 0) ? nC_st1_b165_c0 : nC_st1_b165_c1;
  assign nC_st2_b167_c0 = (nC_st1_b166_c0 == 0) ? nC_st1_b167_c0 : nC_st1_b167_c1;
  assign nC_st2_b169_c0 = (nC_st1_b168_c0 == 0) ? nC_st1_b169_c0 : nC_st1_b169_c1;
  assign nC_st2_b171_c0 = (nC_st1_b170_c0 == 0) ? nC_st1_b171_c0 : nC_st1_b171_c1;
  assign nC_st2_b173_c0 = (nC_st1_b172_c0 == 0) ? nC_st1_b173_c0 : nC_st1_b173_c1;
  assign nC_st2_b175_c0 = (nC_st1_b174_c0 == 0) ? nC_st1_b175_c0 : nC_st1_b175_c1;
  assign nC_st2_b177_c0 = (nC_st1_b176_c0 == 0) ? nC_st1_b177_c0 : nC_st1_b177_c1;
  assign nC_st2_b179_c0 = (nC_st1_b178_c0 == 0) ? nC_st1_b179_c0 : nC_st1_b179_c1;
  assign nC_st2_b181_c0 = (nC_st1_b180_c0 == 0) ? nC_st1_b181_c0 : nC_st1_b181_c1;
  assign nC_st2_b183_c0 = (nC_st1_b182_c0 == 0) ? nC_st1_b183_c0 : nC_st1_b183_c1;
  assign nC_st2_b185_c0 = (nC_st1_b184_c0 == 0) ? nC_st1_b185_c0 : nC_st1_b185_c1;
  assign nC_st2_b187_c0 = (nC_st1_b186_c0 == 0) ? nC_st1_b187_c0 : nC_st1_b187_c1;
  assign nC_st2_b189_c0 = (nC_st1_b188_c0 == 0) ? nC_st1_b189_c0 : nC_st1_b189_c1;
  assign nC_st2_b191_c0 = (nC_st1_b190_c0 == 0) ? nC_st1_b191_c0 : nC_st1_b191_c1;
  assign nC_st2_b193_c0 = (nC_st1_b192_c0 == 0) ? nC_st1_b193_c0 : nC_st1_b193_c1;
  assign nC_st2_b195_c0 = (nC_st1_b194_c0 == 0) ? nC_st1_b195_c0 : nC_st1_b195_c1;
  assign nC_st2_b197_c0 = (nC_st1_b196_c0 == 0) ? nC_st1_b197_c0 : nC_st1_b197_c1;
  assign nC_st2_b199_c0 = (nC_st1_b198_c0 == 0) ? nC_st1_b199_c0 : nC_st1_b199_c1;
  assign nC_st2_b201_c0 = (nC_st1_b200_c0 == 0) ? nC_st1_b201_c0 : nC_st1_b201_c1;
  assign nC_st2_b203_c0 = (nC_st1_b202_c0 == 0) ? nC_st1_b203_c0 : nC_st1_b203_c1;
  assign nC_st2_b205_c0 = (nC_st1_b204_c0 == 0) ? nC_st1_b205_c0 : nC_st1_b205_c1;
  assign nC_st2_b207_c0 = (nC_st1_b206_c0 == 0) ? nC_st1_b207_c0 : nC_st1_b207_c1;
  assign nC_st2_b209_c0 = (nC_st1_b208_c0 == 0) ? nC_st1_b209_c0 : nC_st1_b209_c1;
  assign nC_st2_b211_c0 = (nC_st1_b210_c0 == 0) ? nC_st1_b211_c0 : nC_st1_b211_c1;
  assign nC_st2_b213_c0 = (nC_st1_b212_c0 == 0) ? nC_st1_b213_c0 : nC_st1_b213_c1;
  assign nC_st2_b215_c0 = (nC_st1_b214_c0 == 0) ? nC_st1_b215_c0 : nC_st1_b215_c1;
  assign nC_st2_b217_c0 = (nC_st1_b216_c0 == 0) ? nC_st1_b217_c0 : nC_st1_b217_c1;
  assign nC_st2_b219_c0 = (nC_st1_b218_c0 == 0) ? nC_st1_b219_c0 : nC_st1_b219_c1;
  assign nC_st2_b221_c0 = (nC_st1_b220_c0 == 0) ? nC_st1_b221_c0 : nC_st1_b221_c1;
  assign nC_st2_b223_c0 = (nC_st1_b222_c0 == 0) ? nC_st1_b223_c0 : nC_st1_b223_c1;
  assign nC_st2_b225_c0 = (nC_st1_b224_c0 == 0) ? nC_st1_b225_c0 : nC_st1_b225_c1;
  assign nC_st2_b227_c0 = (nC_st1_b226_c0 == 0) ? nC_st1_b227_c0 : nC_st1_b227_c1;
  assign nC_st2_b229_c0 = (nC_st1_b228_c0 == 0) ? nC_st1_b229_c0 : nC_st1_b229_c1;
  assign nC_st2_b231_c0 = (nC_st1_b230_c0 == 0) ? nC_st1_b231_c0 : nC_st1_b231_c1;
  assign nC_st2_b233_c0 = (nC_st1_b232_c0 == 0) ? nC_st1_b233_c0 : nC_st1_b233_c1;
  assign nC_st2_b235_c0 = (nC_st1_b234_c0 == 0) ? nC_st1_b235_c0 : nC_st1_b235_c1;
  assign nC_st2_b237_c0 = (nC_st1_b236_c0 == 0) ? nC_st1_b237_c0 : nC_st1_b237_c1;
  assign nC_st2_b239_c0 = (nC_st1_b238_c0 == 0) ? nC_st1_b239_c0 : nC_st1_b239_c1;
  assign nC_st2_b241_c0 = (nC_st1_b240_c0 == 0) ? nC_st1_b241_c0 : nC_st1_b241_c1;
  assign nC_st2_b243_c0 = (nC_st1_b242_c0 == 0) ? nC_st1_b243_c0 : nC_st1_b243_c1;
  assign nC_st2_b245_c0 = (nC_st1_b244_c0 == 0) ? nC_st1_b245_c0 : nC_st1_b245_c1;
  assign nC_st2_b247_c0 = (nC_st1_b246_c0 == 0) ? nC_st1_b247_c0 : nC_st1_b247_c1;
  assign nC_st2_b249_c0 = (nC_st1_b248_c0 == 0) ? nC_st1_b249_c0 : nC_st1_b249_c1;
  assign nC_st2_b251_c0 = (nC_st1_b250_c0 == 0) ? nC_st1_b251_c0 : nC_st1_b251_c1;
  assign nC_st2_b253_c0 = (nC_st1_b252_c0 == 0) ? nC_st1_b253_c0 : nC_st1_b253_c1;
  assign nC_st2_b255_c0 = (nC_st1_b254_c0 == 0) ? nC_st1_b255_c0 : nC_st1_b255_c1;
  assign nC_st2_b1_c1 = (nC_st1_b0_c1 == 0) ? nC_st1_b1_c0 : nC_st1_b1_c1;
  assign nC_st2_b3_c1 = (nC_st1_b2_c1 == 0) ? nC_st1_b3_c0 : nC_st1_b3_c1;
  assign nC_st2_b5_c1 = (nC_st1_b4_c1 == 0) ? nC_st1_b5_c0 : nC_st1_b5_c1;
  assign nC_st2_b7_c1 = (nC_st1_b6_c1 == 0) ? nC_st1_b7_c0 : nC_st1_b7_c1;
  assign nC_st2_b9_c1 = (nC_st1_b8_c1 == 0) ? nC_st1_b9_c0 : nC_st1_b9_c1;
  assign nC_st2_b11_c1 = (nC_st1_b10_c1 == 0) ? nC_st1_b11_c0 : nC_st1_b11_c1;
  assign nC_st2_b13_c1 = (nC_st1_b12_c1 == 0) ? nC_st1_b13_c0 : nC_st1_b13_c1;
  assign nC_st2_b15_c1 = (nC_st1_b14_c1 == 0) ? nC_st1_b15_c0 : nC_st1_b15_c1;
  assign nC_st2_b17_c1 = (nC_st1_b16_c1 == 0) ? nC_st1_b17_c0 : nC_st1_b17_c1;
  assign nC_st2_b19_c1 = (nC_st1_b18_c1 == 0) ? nC_st1_b19_c0 : nC_st1_b19_c1;
  assign nC_st2_b21_c1 = (nC_st1_b20_c1 == 0) ? nC_st1_b21_c0 : nC_st1_b21_c1;
  assign nC_st2_b23_c1 = (nC_st1_b22_c1 == 0) ? nC_st1_b23_c0 : nC_st1_b23_c1;
  assign nC_st2_b25_c1 = (nC_st1_b24_c1 == 0) ? nC_st1_b25_c0 : nC_st1_b25_c1;
  assign nC_st2_b27_c1 = (nC_st1_b26_c1 == 0) ? nC_st1_b27_c0 : nC_st1_b27_c1;
  assign nC_st2_b29_c1 = (nC_st1_b28_c1 == 0) ? nC_st1_b29_c0 : nC_st1_b29_c1;
  assign nC_st2_b31_c1 = (nC_st1_b30_c1 == 0) ? nC_st1_b31_c0 : nC_st1_b31_c1;
  assign nC_st2_b33_c1 = (nC_st1_b32_c1 == 0) ? nC_st1_b33_c0 : nC_st1_b33_c1;
  assign nC_st2_b35_c1 = (nC_st1_b34_c1 == 0) ? nC_st1_b35_c0 : nC_st1_b35_c1;
  assign nC_st2_b37_c1 = (nC_st1_b36_c1 == 0) ? nC_st1_b37_c0 : nC_st1_b37_c1;
  assign nC_st2_b39_c1 = (nC_st1_b38_c1 == 0) ? nC_st1_b39_c0 : nC_st1_b39_c1;
  assign nC_st2_b41_c1 = (nC_st1_b40_c1 == 0) ? nC_st1_b41_c0 : nC_st1_b41_c1;
  assign nC_st2_b43_c1 = (nC_st1_b42_c1 == 0) ? nC_st1_b43_c0 : nC_st1_b43_c1;
  assign nC_st2_b45_c1 = (nC_st1_b44_c1 == 0) ? nC_st1_b45_c0 : nC_st1_b45_c1;
  assign nC_st2_b47_c1 = (nC_st1_b46_c1 == 0) ? nC_st1_b47_c0 : nC_st1_b47_c1;
  assign nC_st2_b49_c1 = (nC_st1_b48_c1 == 0) ? nC_st1_b49_c0 : nC_st1_b49_c1;
  assign nC_st2_b51_c1 = (nC_st1_b50_c1 == 0) ? nC_st1_b51_c0 : nC_st1_b51_c1;
  assign nC_st2_b53_c1 = (nC_st1_b52_c1 == 0) ? nC_st1_b53_c0 : nC_st1_b53_c1;
  assign nC_st2_b55_c1 = (nC_st1_b54_c1 == 0) ? nC_st1_b55_c0 : nC_st1_b55_c1;
  assign nC_st2_b57_c1 = (nC_st1_b56_c1 == 0) ? nC_st1_b57_c0 : nC_st1_b57_c1;
  assign nC_st2_b59_c1 = (nC_st1_b58_c1 == 0) ? nC_st1_b59_c0 : nC_st1_b59_c1;
  assign nC_st2_b61_c1 = (nC_st1_b60_c1 == 0) ? nC_st1_b61_c0 : nC_st1_b61_c1;
  assign nC_st2_b63_c1 = (nC_st1_b62_c1 == 0) ? nC_st1_b63_c0 : nC_st1_b63_c1;
  assign nC_st2_b65_c1 = (nC_st1_b64_c1 == 0) ? nC_st1_b65_c0 : nC_st1_b65_c1;
  assign nC_st2_b67_c1 = (nC_st1_b66_c1 == 0) ? nC_st1_b67_c0 : nC_st1_b67_c1;
  assign nC_st2_b69_c1 = (nC_st1_b68_c1 == 0) ? nC_st1_b69_c0 : nC_st1_b69_c1;
  assign nC_st2_b71_c1 = (nC_st1_b70_c1 == 0) ? nC_st1_b71_c0 : nC_st1_b71_c1;
  assign nC_st2_b73_c1 = (nC_st1_b72_c1 == 0) ? nC_st1_b73_c0 : nC_st1_b73_c1;
  assign nC_st2_b75_c1 = (nC_st1_b74_c1 == 0) ? nC_st1_b75_c0 : nC_st1_b75_c1;
  assign nC_st2_b77_c1 = (nC_st1_b76_c1 == 0) ? nC_st1_b77_c0 : nC_st1_b77_c1;
  assign nC_st2_b79_c1 = (nC_st1_b78_c1 == 0) ? nC_st1_b79_c0 : nC_st1_b79_c1;
  assign nC_st2_b81_c1 = (nC_st1_b80_c1 == 0) ? nC_st1_b81_c0 : nC_st1_b81_c1;
  assign nC_st2_b83_c1 = (nC_st1_b82_c1 == 0) ? nC_st1_b83_c0 : nC_st1_b83_c1;
  assign nC_st2_b85_c1 = (nC_st1_b84_c1 == 0) ? nC_st1_b85_c0 : nC_st1_b85_c1;
  assign nC_st2_b87_c1 = (nC_st1_b86_c1 == 0) ? nC_st1_b87_c0 : nC_st1_b87_c1;
  assign nC_st2_b89_c1 = (nC_st1_b88_c1 == 0) ? nC_st1_b89_c0 : nC_st1_b89_c1;
  assign nC_st2_b91_c1 = (nC_st1_b90_c1 == 0) ? nC_st1_b91_c0 : nC_st1_b91_c1;
  assign nC_st2_b93_c1 = (nC_st1_b92_c1 == 0) ? nC_st1_b93_c0 : nC_st1_b93_c1;
  assign nC_st2_b95_c1 = (nC_st1_b94_c1 == 0) ? nC_st1_b95_c0 : nC_st1_b95_c1;
  assign nC_st2_b97_c1 = (nC_st1_b96_c1 == 0) ? nC_st1_b97_c0 : nC_st1_b97_c1;
  assign nC_st2_b99_c1 = (nC_st1_b98_c1 == 0) ? nC_st1_b99_c0 : nC_st1_b99_c1;
  assign nC_st2_b101_c1 = (nC_st1_b100_c1 == 0) ? nC_st1_b101_c0 : nC_st1_b101_c1;
  assign nC_st2_b103_c1 = (nC_st1_b102_c1 == 0) ? nC_st1_b103_c0 : nC_st1_b103_c1;
  assign nC_st2_b105_c1 = (nC_st1_b104_c1 == 0) ? nC_st1_b105_c0 : nC_st1_b105_c1;
  assign nC_st2_b107_c1 = (nC_st1_b106_c1 == 0) ? nC_st1_b107_c0 : nC_st1_b107_c1;
  assign nC_st2_b109_c1 = (nC_st1_b108_c1 == 0) ? nC_st1_b109_c0 : nC_st1_b109_c1;
  assign nC_st2_b111_c1 = (nC_st1_b110_c1 == 0) ? nC_st1_b111_c0 : nC_st1_b111_c1;
  assign nC_st2_b113_c1 = (nC_st1_b112_c1 == 0) ? nC_st1_b113_c0 : nC_st1_b113_c1;
  assign nC_st2_b115_c1 = (nC_st1_b114_c1 == 0) ? nC_st1_b115_c0 : nC_st1_b115_c1;
  assign nC_st2_b117_c1 = (nC_st1_b116_c1 == 0) ? nC_st1_b117_c0 : nC_st1_b117_c1;
  assign nC_st2_b119_c1 = (nC_st1_b118_c1 == 0) ? nC_st1_b119_c0 : nC_st1_b119_c1;
  assign nC_st2_b121_c1 = (nC_st1_b120_c1 == 0) ? nC_st1_b121_c0 : nC_st1_b121_c1;
  assign nC_st2_b123_c1 = (nC_st1_b122_c1 == 0) ? nC_st1_b123_c0 : nC_st1_b123_c1;
  assign nC_st2_b125_c1 = (nC_st1_b124_c1 == 0) ? nC_st1_b125_c0 : nC_st1_b125_c1;
  assign nC_st2_b127_c1 = (nC_st1_b126_c1 == 0) ? nC_st1_b127_c0 : nC_st1_b127_c1;
  assign nC_st2_b129_c1 = (nC_st1_b128_c1 == 0) ? nC_st1_b129_c0 : nC_st1_b129_c1;
  assign nC_st2_b131_c1 = (nC_st1_b130_c1 == 0) ? nC_st1_b131_c0 : nC_st1_b131_c1;
  assign nC_st2_b133_c1 = (nC_st1_b132_c1 == 0) ? nC_st1_b133_c0 : nC_st1_b133_c1;
  assign nC_st2_b135_c1 = (nC_st1_b134_c1 == 0) ? nC_st1_b135_c0 : nC_st1_b135_c1;
  assign nC_st2_b137_c1 = (nC_st1_b136_c1 == 0) ? nC_st1_b137_c0 : nC_st1_b137_c1;
  assign nC_st2_b139_c1 = (nC_st1_b138_c1 == 0) ? nC_st1_b139_c0 : nC_st1_b139_c1;
  assign nC_st2_b141_c1 = (nC_st1_b140_c1 == 0) ? nC_st1_b141_c0 : nC_st1_b141_c1;
  assign nC_st2_b143_c1 = (nC_st1_b142_c1 == 0) ? nC_st1_b143_c0 : nC_st1_b143_c1;
  assign nC_st2_b145_c1 = (nC_st1_b144_c1 == 0) ? nC_st1_b145_c0 : nC_st1_b145_c1;
  assign nC_st2_b147_c1 = (nC_st1_b146_c1 == 0) ? nC_st1_b147_c0 : nC_st1_b147_c1;
  assign nC_st2_b149_c1 = (nC_st1_b148_c1 == 0) ? nC_st1_b149_c0 : nC_st1_b149_c1;
  assign nC_st2_b151_c1 = (nC_st1_b150_c1 == 0) ? nC_st1_b151_c0 : nC_st1_b151_c1;
  assign nC_st2_b153_c1 = (nC_st1_b152_c1 == 0) ? nC_st1_b153_c0 : nC_st1_b153_c1;
  assign nC_st2_b155_c1 = (nC_st1_b154_c1 == 0) ? nC_st1_b155_c0 : nC_st1_b155_c1;
  assign nC_st2_b157_c1 = (nC_st1_b156_c1 == 0) ? nC_st1_b157_c0 : nC_st1_b157_c1;
  assign nC_st2_b159_c1 = (nC_st1_b158_c1 == 0) ? nC_st1_b159_c0 : nC_st1_b159_c1;
  assign nC_st2_b161_c1 = (nC_st1_b160_c1 == 0) ? nC_st1_b161_c0 : nC_st1_b161_c1;
  assign nC_st2_b163_c1 = (nC_st1_b162_c1 == 0) ? nC_st1_b163_c0 : nC_st1_b163_c1;
  assign nC_st2_b165_c1 = (nC_st1_b164_c1 == 0) ? nC_st1_b165_c0 : nC_st1_b165_c1;
  assign nC_st2_b167_c1 = (nC_st1_b166_c1 == 0) ? nC_st1_b167_c0 : nC_st1_b167_c1;
  assign nC_st2_b169_c1 = (nC_st1_b168_c1 == 0) ? nC_st1_b169_c0 : nC_st1_b169_c1;
  assign nC_st2_b171_c1 = (nC_st1_b170_c1 == 0) ? nC_st1_b171_c0 : nC_st1_b171_c1;
  assign nC_st2_b173_c1 = (nC_st1_b172_c1 == 0) ? nC_st1_b173_c0 : nC_st1_b173_c1;
  assign nC_st2_b175_c1 = (nC_st1_b174_c1 == 0) ? nC_st1_b175_c0 : nC_st1_b175_c1;
  assign nC_st2_b177_c1 = (nC_st1_b176_c1 == 0) ? nC_st1_b177_c0 : nC_st1_b177_c1;
  assign nC_st2_b179_c1 = (nC_st1_b178_c1 == 0) ? nC_st1_b179_c0 : nC_st1_b179_c1;
  assign nC_st2_b181_c1 = (nC_st1_b180_c1 == 0) ? nC_st1_b181_c0 : nC_st1_b181_c1;
  assign nC_st2_b183_c1 = (nC_st1_b182_c1 == 0) ? nC_st1_b183_c0 : nC_st1_b183_c1;
  assign nC_st2_b185_c1 = (nC_st1_b184_c1 == 0) ? nC_st1_b185_c0 : nC_st1_b185_c1;
  assign nC_st2_b187_c1 = (nC_st1_b186_c1 == 0) ? nC_st1_b187_c0 : nC_st1_b187_c1;
  assign nC_st2_b189_c1 = (nC_st1_b188_c1 == 0) ? nC_st1_b189_c0 : nC_st1_b189_c1;
  assign nC_st2_b191_c1 = (nC_st1_b190_c1 == 0) ? nC_st1_b191_c0 : nC_st1_b191_c1;
  assign nC_st2_b193_c1 = (nC_st1_b192_c1 == 0) ? nC_st1_b193_c0 : nC_st1_b193_c1;
  assign nC_st2_b195_c1 = (nC_st1_b194_c1 == 0) ? nC_st1_b195_c0 : nC_st1_b195_c1;
  assign nC_st2_b197_c1 = (nC_st1_b196_c1 == 0) ? nC_st1_b197_c0 : nC_st1_b197_c1;
  assign nC_st2_b199_c1 = (nC_st1_b198_c1 == 0) ? nC_st1_b199_c0 : nC_st1_b199_c1;
  assign nC_st2_b201_c1 = (nC_st1_b200_c1 == 0) ? nC_st1_b201_c0 : nC_st1_b201_c1;
  assign nC_st2_b203_c1 = (nC_st1_b202_c1 == 0) ? nC_st1_b203_c0 : nC_st1_b203_c1;
  assign nC_st2_b205_c1 = (nC_st1_b204_c1 == 0) ? nC_st1_b205_c0 : nC_st1_b205_c1;
  assign nC_st2_b207_c1 = (nC_st1_b206_c1 == 0) ? nC_st1_b207_c0 : nC_st1_b207_c1;
  assign nC_st2_b209_c1 = (nC_st1_b208_c1 == 0) ? nC_st1_b209_c0 : nC_st1_b209_c1;
  assign nC_st2_b211_c1 = (nC_st1_b210_c1 == 0) ? nC_st1_b211_c0 : nC_st1_b211_c1;
  assign nC_st2_b213_c1 = (nC_st1_b212_c1 == 0) ? nC_st1_b213_c0 : nC_st1_b213_c1;
  assign nC_st2_b215_c1 = (nC_st1_b214_c1 == 0) ? nC_st1_b215_c0 : nC_st1_b215_c1;
  assign nC_st2_b217_c1 = (nC_st1_b216_c1 == 0) ? nC_st1_b217_c0 : nC_st1_b217_c1;
  assign nC_st2_b219_c1 = (nC_st1_b218_c1 == 0) ? nC_st1_b219_c0 : nC_st1_b219_c1;
  assign nC_st2_b221_c1 = (nC_st1_b220_c1 == 0) ? nC_st1_b221_c0 : nC_st1_b221_c1;
  assign nC_st2_b223_c1 = (nC_st1_b222_c1 == 0) ? nC_st1_b223_c0 : nC_st1_b223_c1;
  assign nC_st2_b225_c1 = (nC_st1_b224_c1 == 0) ? nC_st1_b225_c0 : nC_st1_b225_c1;
  assign nC_st2_b227_c1 = (nC_st1_b226_c1 == 0) ? nC_st1_b227_c0 : nC_st1_b227_c1;
  assign nC_st2_b229_c1 = (nC_st1_b228_c1 == 0) ? nC_st1_b229_c0 : nC_st1_b229_c1;
  assign nC_st2_b231_c1 = (nC_st1_b230_c1 == 0) ? nC_st1_b231_c0 : nC_st1_b231_c1;
  assign nC_st2_b233_c1 = (nC_st1_b232_c1 == 0) ? nC_st1_b233_c0 : nC_st1_b233_c1;
  assign nC_st2_b235_c1 = (nC_st1_b234_c1 == 0) ? nC_st1_b235_c0 : nC_st1_b235_c1;
  assign nC_st2_b237_c1 = (nC_st1_b236_c1 == 0) ? nC_st1_b237_c0 : nC_st1_b237_c1;
  assign nC_st2_b239_c1 = (nC_st1_b238_c1 == 0) ? nC_st1_b239_c0 : nC_st1_b239_c1;
  assign nC_st2_b241_c1 = (nC_st1_b240_c1 == 0) ? nC_st1_b241_c0 : nC_st1_b241_c1;
  assign nC_st2_b243_c1 = (nC_st1_b242_c1 == 0) ? nC_st1_b243_c0 : nC_st1_b243_c1;
  assign nC_st2_b245_c1 = (nC_st1_b244_c1 == 0) ? nC_st1_b245_c0 : nC_st1_b245_c1;
  assign nC_st2_b247_c1 = (nC_st1_b246_c1 == 0) ? nC_st1_b247_c0 : nC_st1_b247_c1;
  assign nC_st2_b249_c1 = (nC_st1_b248_c1 == 0) ? nC_st1_b249_c0 : nC_st1_b249_c1;
  assign nC_st2_b251_c1 = (nC_st1_b250_c1 == 0) ? nC_st1_b251_c0 : nC_st1_b251_c1;
  assign nC_st2_b253_c1 = (nC_st1_b252_c1 == 0) ? nC_st1_b253_c0 : nC_st1_b253_c1;
  assign nC_st2_b255_c1 = (nC_st1_b254_c1 == 0) ? nC_st1_b255_c0 : nC_st1_b255_c1;

  assign nS_st3_b0_c0 = nS_st2_b0_c0;
  assign nS_st3_b1_c0 = nS_st2_b1_c0;
  assign nS_st3_b2_c0 = (nC_st2_b1_c0 == 0) ? nS_st2_b2_c0 : nS_st2_b2_c1;
  assign nS_st3_b3_c0 = (nC_st2_b1_c0 == 0) ? nS_st2_b3_c0 : nS_st2_b3_c1;
  assign nS_st3_b4_c0 = nS_st2_b4_c0;
  assign nS_st3_b5_c0 = nS_st2_b5_c0;
  assign nS_st3_b6_c0 = (nC_st2_b5_c0 == 0) ? nS_st2_b6_c0 : nS_st2_b6_c1;
  assign nS_st3_b7_c0 = (nC_st2_b5_c0 == 0) ? nS_st2_b7_c0 : nS_st2_b7_c1;
  assign nS_st3_b8_c0 = nS_st2_b8_c0;
  assign nS_st3_b9_c0 = nS_st2_b9_c0;
  assign nS_st3_b10_c0 = (nC_st2_b9_c0 == 0) ? nS_st2_b10_c0 : nS_st2_b10_c1;
  assign nS_st3_b11_c0 = (nC_st2_b9_c0 == 0) ? nS_st2_b11_c0 : nS_st2_b11_c1;
  assign nS_st3_b12_c0 = nS_st2_b12_c0;
  assign nS_st3_b13_c0 = nS_st2_b13_c0;
  assign nS_st3_b14_c0 = (nC_st2_b13_c0 == 0) ? nS_st2_b14_c0 : nS_st2_b14_c1;
  assign nS_st3_b15_c0 = (nC_st2_b13_c0 == 0) ? nS_st2_b15_c0 : nS_st2_b15_c1;
  assign nS_st3_b16_c0 = nS_st2_b16_c0;
  assign nS_st3_b17_c0 = nS_st2_b17_c0;
  assign nS_st3_b18_c0 = (nC_st2_b17_c0 == 0) ? nS_st2_b18_c0 : nS_st2_b18_c1;
  assign nS_st3_b19_c0 = (nC_st2_b17_c0 == 0) ? nS_st2_b19_c0 : nS_st2_b19_c1;
  assign nS_st3_b20_c0 = nS_st2_b20_c0;
  assign nS_st3_b21_c0 = nS_st2_b21_c0;
  assign nS_st3_b22_c0 = (nC_st2_b21_c0 == 0) ? nS_st2_b22_c0 : nS_st2_b22_c1;
  assign nS_st3_b23_c0 = (nC_st2_b21_c0 == 0) ? nS_st2_b23_c0 : nS_st2_b23_c1;
  assign nS_st3_b24_c0 = nS_st2_b24_c0;
  assign nS_st3_b25_c0 = nS_st2_b25_c0;
  assign nS_st3_b26_c0 = (nC_st2_b25_c0 == 0) ? nS_st2_b26_c0 : nS_st2_b26_c1;
  assign nS_st3_b27_c0 = (nC_st2_b25_c0 == 0) ? nS_st2_b27_c0 : nS_st2_b27_c1;
  assign nS_st3_b28_c0 = nS_st2_b28_c0;
  assign nS_st3_b29_c0 = nS_st2_b29_c0;
  assign nS_st3_b30_c0 = (nC_st2_b29_c0 == 0) ? nS_st2_b30_c0 : nS_st2_b30_c1;
  assign nS_st3_b31_c0 = (nC_st2_b29_c0 == 0) ? nS_st2_b31_c0 : nS_st2_b31_c1;
  assign nS_st3_b32_c0 = nS_st2_b32_c0;
  assign nS_st3_b33_c0 = nS_st2_b33_c0;
  assign nS_st3_b34_c0 = (nC_st2_b33_c0 == 0) ? nS_st2_b34_c0 : nS_st2_b34_c1;
  assign nS_st3_b35_c0 = (nC_st2_b33_c0 == 0) ? nS_st2_b35_c0 : nS_st2_b35_c1;
  assign nS_st3_b36_c0 = nS_st2_b36_c0;
  assign nS_st3_b37_c0 = nS_st2_b37_c0;
  assign nS_st3_b38_c0 = (nC_st2_b37_c0 == 0) ? nS_st2_b38_c0 : nS_st2_b38_c1;
  assign nS_st3_b39_c0 = (nC_st2_b37_c0 == 0) ? nS_st2_b39_c0 : nS_st2_b39_c1;
  assign nS_st3_b40_c0 = nS_st2_b40_c0;
  assign nS_st3_b41_c0 = nS_st2_b41_c0;
  assign nS_st3_b42_c0 = (nC_st2_b41_c0 == 0) ? nS_st2_b42_c0 : nS_st2_b42_c1;
  assign nS_st3_b43_c0 = (nC_st2_b41_c0 == 0) ? nS_st2_b43_c0 : nS_st2_b43_c1;
  assign nS_st3_b44_c0 = nS_st2_b44_c0;
  assign nS_st3_b45_c0 = nS_st2_b45_c0;
  assign nS_st3_b46_c0 = (nC_st2_b45_c0 == 0) ? nS_st2_b46_c0 : nS_st2_b46_c1;
  assign nS_st3_b47_c0 = (nC_st2_b45_c0 == 0) ? nS_st2_b47_c0 : nS_st2_b47_c1;
  assign nS_st3_b48_c0 = nS_st2_b48_c0;
  assign nS_st3_b49_c0 = nS_st2_b49_c0;
  assign nS_st3_b50_c0 = (nC_st2_b49_c0 == 0) ? nS_st2_b50_c0 : nS_st2_b50_c1;
  assign nS_st3_b51_c0 = (nC_st2_b49_c0 == 0) ? nS_st2_b51_c0 : nS_st2_b51_c1;
  assign nS_st3_b52_c0 = nS_st2_b52_c0;
  assign nS_st3_b53_c0 = nS_st2_b53_c0;
  assign nS_st3_b54_c0 = (nC_st2_b53_c0 == 0) ? nS_st2_b54_c0 : nS_st2_b54_c1;
  assign nS_st3_b55_c0 = (nC_st2_b53_c0 == 0) ? nS_st2_b55_c0 : nS_st2_b55_c1;
  assign nS_st3_b56_c0 = nS_st2_b56_c0;
  assign nS_st3_b57_c0 = nS_st2_b57_c0;
  assign nS_st3_b58_c0 = (nC_st2_b57_c0 == 0) ? nS_st2_b58_c0 : nS_st2_b58_c1;
  assign nS_st3_b59_c0 = (nC_st2_b57_c0 == 0) ? nS_st2_b59_c0 : nS_st2_b59_c1;
  assign nS_st3_b60_c0 = nS_st2_b60_c0;
  assign nS_st3_b61_c0 = nS_st2_b61_c0;
  assign nS_st3_b62_c0 = (nC_st2_b61_c0 == 0) ? nS_st2_b62_c0 : nS_st2_b62_c1;
  assign nS_st3_b63_c0 = (nC_st2_b61_c0 == 0) ? nS_st2_b63_c0 : nS_st2_b63_c1;
  assign nS_st3_b64_c0 = nS_st2_b64_c0;
  assign nS_st3_b65_c0 = nS_st2_b65_c0;
  assign nS_st3_b66_c0 = (nC_st2_b65_c0 == 0) ? nS_st2_b66_c0 : nS_st2_b66_c1;
  assign nS_st3_b67_c0 = (nC_st2_b65_c0 == 0) ? nS_st2_b67_c0 : nS_st2_b67_c1;
  assign nS_st3_b68_c0 = nS_st2_b68_c0;
  assign nS_st3_b69_c0 = nS_st2_b69_c0;
  assign nS_st3_b70_c0 = (nC_st2_b69_c0 == 0) ? nS_st2_b70_c0 : nS_st2_b70_c1;
  assign nS_st3_b71_c0 = (nC_st2_b69_c0 == 0) ? nS_st2_b71_c0 : nS_st2_b71_c1;
  assign nS_st3_b72_c0 = nS_st2_b72_c0;
  assign nS_st3_b73_c0 = nS_st2_b73_c0;
  assign nS_st3_b74_c0 = (nC_st2_b73_c0 == 0) ? nS_st2_b74_c0 : nS_st2_b74_c1;
  assign nS_st3_b75_c0 = (nC_st2_b73_c0 == 0) ? nS_st2_b75_c0 : nS_st2_b75_c1;
  assign nS_st3_b76_c0 = nS_st2_b76_c0;
  assign nS_st3_b77_c0 = nS_st2_b77_c0;
  assign nS_st3_b78_c0 = (nC_st2_b77_c0 == 0) ? nS_st2_b78_c0 : nS_st2_b78_c1;
  assign nS_st3_b79_c0 = (nC_st2_b77_c0 == 0) ? nS_st2_b79_c0 : nS_st2_b79_c1;
  assign nS_st3_b80_c0 = nS_st2_b80_c0;
  assign nS_st3_b81_c0 = nS_st2_b81_c0;
  assign nS_st3_b82_c0 = (nC_st2_b81_c0 == 0) ? nS_st2_b82_c0 : nS_st2_b82_c1;
  assign nS_st3_b83_c0 = (nC_st2_b81_c0 == 0) ? nS_st2_b83_c0 : nS_st2_b83_c1;
  assign nS_st3_b84_c0 = nS_st2_b84_c0;
  assign nS_st3_b85_c0 = nS_st2_b85_c0;
  assign nS_st3_b86_c0 = (nC_st2_b85_c0 == 0) ? nS_st2_b86_c0 : nS_st2_b86_c1;
  assign nS_st3_b87_c0 = (nC_st2_b85_c0 == 0) ? nS_st2_b87_c0 : nS_st2_b87_c1;
  assign nS_st3_b88_c0 = nS_st2_b88_c0;
  assign nS_st3_b89_c0 = nS_st2_b89_c0;
  assign nS_st3_b90_c0 = (nC_st2_b89_c0 == 0) ? nS_st2_b90_c0 : nS_st2_b90_c1;
  assign nS_st3_b91_c0 = (nC_st2_b89_c0 == 0) ? nS_st2_b91_c0 : nS_st2_b91_c1;
  assign nS_st3_b92_c0 = nS_st2_b92_c0;
  assign nS_st3_b93_c0 = nS_st2_b93_c0;
  assign nS_st3_b94_c0 = (nC_st2_b93_c0 == 0) ? nS_st2_b94_c0 : nS_st2_b94_c1;
  assign nS_st3_b95_c0 = (nC_st2_b93_c0 == 0) ? nS_st2_b95_c0 : nS_st2_b95_c1;
  assign nS_st3_b96_c0 = nS_st2_b96_c0;
  assign nS_st3_b97_c0 = nS_st2_b97_c0;
  assign nS_st3_b98_c0 = (nC_st2_b97_c0 == 0) ? nS_st2_b98_c0 : nS_st2_b98_c1;
  assign nS_st3_b99_c0 = (nC_st2_b97_c0 == 0) ? nS_st2_b99_c0 : nS_st2_b99_c1;
  assign nS_st3_b100_c0 = nS_st2_b100_c0;
  assign nS_st3_b101_c0 = nS_st2_b101_c0;
  assign nS_st3_b102_c0 = (nC_st2_b101_c0 == 0) ? nS_st2_b102_c0 : nS_st2_b102_c1;
  assign nS_st3_b103_c0 = (nC_st2_b101_c0 == 0) ? nS_st2_b103_c0 : nS_st2_b103_c1;
  assign nS_st3_b104_c0 = nS_st2_b104_c0;
  assign nS_st3_b105_c0 = nS_st2_b105_c0;
  assign nS_st3_b106_c0 = (nC_st2_b105_c0 == 0) ? nS_st2_b106_c0 : nS_st2_b106_c1;
  assign nS_st3_b107_c0 = (nC_st2_b105_c0 == 0) ? nS_st2_b107_c0 : nS_st2_b107_c1;
  assign nS_st3_b108_c0 = nS_st2_b108_c0;
  assign nS_st3_b109_c0 = nS_st2_b109_c0;
  assign nS_st3_b110_c0 = (nC_st2_b109_c0 == 0) ? nS_st2_b110_c0 : nS_st2_b110_c1;
  assign nS_st3_b111_c0 = (nC_st2_b109_c0 == 0) ? nS_st2_b111_c0 : nS_st2_b111_c1;
  assign nS_st3_b112_c0 = nS_st2_b112_c0;
  assign nS_st3_b113_c0 = nS_st2_b113_c0;
  assign nS_st3_b114_c0 = (nC_st2_b113_c0 == 0) ? nS_st2_b114_c0 : nS_st2_b114_c1;
  assign nS_st3_b115_c0 = (nC_st2_b113_c0 == 0) ? nS_st2_b115_c0 : nS_st2_b115_c1;
  assign nS_st3_b116_c0 = nS_st2_b116_c0;
  assign nS_st3_b117_c0 = nS_st2_b117_c0;
  assign nS_st3_b118_c0 = (nC_st2_b117_c0 == 0) ? nS_st2_b118_c0 : nS_st2_b118_c1;
  assign nS_st3_b119_c0 = (nC_st2_b117_c0 == 0) ? nS_st2_b119_c0 : nS_st2_b119_c1;
  assign nS_st3_b120_c0 = nS_st2_b120_c0;
  assign nS_st3_b121_c0 = nS_st2_b121_c0;
  assign nS_st3_b122_c0 = (nC_st2_b121_c0 == 0) ? nS_st2_b122_c0 : nS_st2_b122_c1;
  assign nS_st3_b123_c0 = (nC_st2_b121_c0 == 0) ? nS_st2_b123_c0 : nS_st2_b123_c1;
  assign nS_st3_b124_c0 = nS_st2_b124_c0;
  assign nS_st3_b125_c0 = nS_st2_b125_c0;
  assign nS_st3_b126_c0 = (nC_st2_b125_c0 == 0) ? nS_st2_b126_c0 : nS_st2_b126_c1;
  assign nS_st3_b127_c0 = (nC_st2_b125_c0 == 0) ? nS_st2_b127_c0 : nS_st2_b127_c1;
  assign nS_st3_b128_c0 = nS_st2_b128_c0;
  assign nS_st3_b129_c0 = nS_st2_b129_c0;
  assign nS_st3_b130_c0 = (nC_st2_b129_c0 == 0) ? nS_st2_b130_c0 : nS_st2_b130_c1;
  assign nS_st3_b131_c0 = (nC_st2_b129_c0 == 0) ? nS_st2_b131_c0 : nS_st2_b131_c1;
  assign nS_st3_b132_c0 = nS_st2_b132_c0;
  assign nS_st3_b133_c0 = nS_st2_b133_c0;
  assign nS_st3_b134_c0 = (nC_st2_b133_c0 == 0) ? nS_st2_b134_c0 : nS_st2_b134_c1;
  assign nS_st3_b135_c0 = (nC_st2_b133_c0 == 0) ? nS_st2_b135_c0 : nS_st2_b135_c1;
  assign nS_st3_b136_c0 = nS_st2_b136_c0;
  assign nS_st3_b137_c0 = nS_st2_b137_c0;
  assign nS_st3_b138_c0 = (nC_st2_b137_c0 == 0) ? nS_st2_b138_c0 : nS_st2_b138_c1;
  assign nS_st3_b139_c0 = (nC_st2_b137_c0 == 0) ? nS_st2_b139_c0 : nS_st2_b139_c1;
  assign nS_st3_b140_c0 = nS_st2_b140_c0;
  assign nS_st3_b141_c0 = nS_st2_b141_c0;
  assign nS_st3_b142_c0 = (nC_st2_b141_c0 == 0) ? nS_st2_b142_c0 : nS_st2_b142_c1;
  assign nS_st3_b143_c0 = (nC_st2_b141_c0 == 0) ? nS_st2_b143_c0 : nS_st2_b143_c1;
  assign nS_st3_b144_c0 = nS_st2_b144_c0;
  assign nS_st3_b145_c0 = nS_st2_b145_c0;
  assign nS_st3_b146_c0 = (nC_st2_b145_c0 == 0) ? nS_st2_b146_c0 : nS_st2_b146_c1;
  assign nS_st3_b147_c0 = (nC_st2_b145_c0 == 0) ? nS_st2_b147_c0 : nS_st2_b147_c1;
  assign nS_st3_b148_c0 = nS_st2_b148_c0;
  assign nS_st3_b149_c0 = nS_st2_b149_c0;
  assign nS_st3_b150_c0 = (nC_st2_b149_c0 == 0) ? nS_st2_b150_c0 : nS_st2_b150_c1;
  assign nS_st3_b151_c0 = (nC_st2_b149_c0 == 0) ? nS_st2_b151_c0 : nS_st2_b151_c1;
  assign nS_st3_b152_c0 = nS_st2_b152_c0;
  assign nS_st3_b153_c0 = nS_st2_b153_c0;
  assign nS_st3_b154_c0 = (nC_st2_b153_c0 == 0) ? nS_st2_b154_c0 : nS_st2_b154_c1;
  assign nS_st3_b155_c0 = (nC_st2_b153_c0 == 0) ? nS_st2_b155_c0 : nS_st2_b155_c1;
  assign nS_st3_b156_c0 = nS_st2_b156_c0;
  assign nS_st3_b157_c0 = nS_st2_b157_c0;
  assign nS_st3_b158_c0 = (nC_st2_b157_c0 == 0) ? nS_st2_b158_c0 : nS_st2_b158_c1;
  assign nS_st3_b159_c0 = (nC_st2_b157_c0 == 0) ? nS_st2_b159_c0 : nS_st2_b159_c1;
  assign nS_st3_b160_c0 = nS_st2_b160_c0;
  assign nS_st3_b161_c0 = nS_st2_b161_c0;
  assign nS_st3_b162_c0 = (nC_st2_b161_c0 == 0) ? nS_st2_b162_c0 : nS_st2_b162_c1;
  assign nS_st3_b163_c0 = (nC_st2_b161_c0 == 0) ? nS_st2_b163_c0 : nS_st2_b163_c1;
  assign nS_st3_b164_c0 = nS_st2_b164_c0;
  assign nS_st3_b165_c0 = nS_st2_b165_c0;
  assign nS_st3_b166_c0 = (nC_st2_b165_c0 == 0) ? nS_st2_b166_c0 : nS_st2_b166_c1;
  assign nS_st3_b167_c0 = (nC_st2_b165_c0 == 0) ? nS_st2_b167_c0 : nS_st2_b167_c1;
  assign nS_st3_b168_c0 = nS_st2_b168_c0;
  assign nS_st3_b169_c0 = nS_st2_b169_c0;
  assign nS_st3_b170_c0 = (nC_st2_b169_c0 == 0) ? nS_st2_b170_c0 : nS_st2_b170_c1;
  assign nS_st3_b171_c0 = (nC_st2_b169_c0 == 0) ? nS_st2_b171_c0 : nS_st2_b171_c1;
  assign nS_st3_b172_c0 = nS_st2_b172_c0;
  assign nS_st3_b173_c0 = nS_st2_b173_c0;
  assign nS_st3_b174_c0 = (nC_st2_b173_c0 == 0) ? nS_st2_b174_c0 : nS_st2_b174_c1;
  assign nS_st3_b175_c0 = (nC_st2_b173_c0 == 0) ? nS_st2_b175_c0 : nS_st2_b175_c1;
  assign nS_st3_b176_c0 = nS_st2_b176_c0;
  assign nS_st3_b177_c0 = nS_st2_b177_c0;
  assign nS_st3_b178_c0 = (nC_st2_b177_c0 == 0) ? nS_st2_b178_c0 : nS_st2_b178_c1;
  assign nS_st3_b179_c0 = (nC_st2_b177_c0 == 0) ? nS_st2_b179_c0 : nS_st2_b179_c1;
  assign nS_st3_b180_c0 = nS_st2_b180_c0;
  assign nS_st3_b181_c0 = nS_st2_b181_c0;
  assign nS_st3_b182_c0 = (nC_st2_b181_c0 == 0) ? nS_st2_b182_c0 : nS_st2_b182_c1;
  assign nS_st3_b183_c0 = (nC_st2_b181_c0 == 0) ? nS_st2_b183_c0 : nS_st2_b183_c1;
  assign nS_st3_b184_c0 = nS_st2_b184_c0;
  assign nS_st3_b185_c0 = nS_st2_b185_c0;
  assign nS_st3_b186_c0 = (nC_st2_b185_c0 == 0) ? nS_st2_b186_c0 : nS_st2_b186_c1;
  assign nS_st3_b187_c0 = (nC_st2_b185_c0 == 0) ? nS_st2_b187_c0 : nS_st2_b187_c1;
  assign nS_st3_b188_c0 = nS_st2_b188_c0;
  assign nS_st3_b189_c0 = nS_st2_b189_c0;
  assign nS_st3_b190_c0 = (nC_st2_b189_c0 == 0) ? nS_st2_b190_c0 : nS_st2_b190_c1;
  assign nS_st3_b191_c0 = (nC_st2_b189_c0 == 0) ? nS_st2_b191_c0 : nS_st2_b191_c1;
  assign nS_st3_b192_c0 = nS_st2_b192_c0;
  assign nS_st3_b193_c0 = nS_st2_b193_c0;
  assign nS_st3_b194_c0 = (nC_st2_b193_c0 == 0) ? nS_st2_b194_c0 : nS_st2_b194_c1;
  assign nS_st3_b195_c0 = (nC_st2_b193_c0 == 0) ? nS_st2_b195_c0 : nS_st2_b195_c1;
  assign nS_st3_b196_c0 = nS_st2_b196_c0;
  assign nS_st3_b197_c0 = nS_st2_b197_c0;
  assign nS_st3_b198_c0 = (nC_st2_b197_c0 == 0) ? nS_st2_b198_c0 : nS_st2_b198_c1;
  assign nS_st3_b199_c0 = (nC_st2_b197_c0 == 0) ? nS_st2_b199_c0 : nS_st2_b199_c1;
  assign nS_st3_b200_c0 = nS_st2_b200_c0;
  assign nS_st3_b201_c0 = nS_st2_b201_c0;
  assign nS_st3_b202_c0 = (nC_st2_b201_c0 == 0) ? nS_st2_b202_c0 : nS_st2_b202_c1;
  assign nS_st3_b203_c0 = (nC_st2_b201_c0 == 0) ? nS_st2_b203_c0 : nS_st2_b203_c1;
  assign nS_st3_b204_c0 = nS_st2_b204_c0;
  assign nS_st3_b205_c0 = nS_st2_b205_c0;
  assign nS_st3_b206_c0 = (nC_st2_b205_c0 == 0) ? nS_st2_b206_c0 : nS_st2_b206_c1;
  assign nS_st3_b207_c0 = (nC_st2_b205_c0 == 0) ? nS_st2_b207_c0 : nS_st2_b207_c1;
  assign nS_st3_b208_c0 = nS_st2_b208_c0;
  assign nS_st3_b209_c0 = nS_st2_b209_c0;
  assign nS_st3_b210_c0 = (nC_st2_b209_c0 == 0) ? nS_st2_b210_c0 : nS_st2_b210_c1;
  assign nS_st3_b211_c0 = (nC_st2_b209_c0 == 0) ? nS_st2_b211_c0 : nS_st2_b211_c1;
  assign nS_st3_b212_c0 = nS_st2_b212_c0;
  assign nS_st3_b213_c0 = nS_st2_b213_c0;
  assign nS_st3_b214_c0 = (nC_st2_b213_c0 == 0) ? nS_st2_b214_c0 : nS_st2_b214_c1;
  assign nS_st3_b215_c0 = (nC_st2_b213_c0 == 0) ? nS_st2_b215_c0 : nS_st2_b215_c1;
  assign nS_st3_b216_c0 = nS_st2_b216_c0;
  assign nS_st3_b217_c0 = nS_st2_b217_c0;
  assign nS_st3_b218_c0 = (nC_st2_b217_c0 == 0) ? nS_st2_b218_c0 : nS_st2_b218_c1;
  assign nS_st3_b219_c0 = (nC_st2_b217_c0 == 0) ? nS_st2_b219_c0 : nS_st2_b219_c1;
  assign nS_st3_b220_c0 = nS_st2_b220_c0;
  assign nS_st3_b221_c0 = nS_st2_b221_c0;
  assign nS_st3_b222_c0 = (nC_st2_b221_c0 == 0) ? nS_st2_b222_c0 : nS_st2_b222_c1;
  assign nS_st3_b223_c0 = (nC_st2_b221_c0 == 0) ? nS_st2_b223_c0 : nS_st2_b223_c1;
  assign nS_st3_b224_c0 = nS_st2_b224_c0;
  assign nS_st3_b225_c0 = nS_st2_b225_c0;
  assign nS_st3_b226_c0 = (nC_st2_b225_c0 == 0) ? nS_st2_b226_c0 : nS_st2_b226_c1;
  assign nS_st3_b227_c0 = (nC_st2_b225_c0 == 0) ? nS_st2_b227_c0 : nS_st2_b227_c1;
  assign nS_st3_b228_c0 = nS_st2_b228_c0;
  assign nS_st3_b229_c0 = nS_st2_b229_c0;
  assign nS_st3_b230_c0 = (nC_st2_b229_c0 == 0) ? nS_st2_b230_c0 : nS_st2_b230_c1;
  assign nS_st3_b231_c0 = (nC_st2_b229_c0 == 0) ? nS_st2_b231_c0 : nS_st2_b231_c1;
  assign nS_st3_b232_c0 = nS_st2_b232_c0;
  assign nS_st3_b233_c0 = nS_st2_b233_c0;
  assign nS_st3_b234_c0 = (nC_st2_b233_c0 == 0) ? nS_st2_b234_c0 : nS_st2_b234_c1;
  assign nS_st3_b235_c0 = (nC_st2_b233_c0 == 0) ? nS_st2_b235_c0 : nS_st2_b235_c1;
  assign nS_st3_b236_c0 = nS_st2_b236_c0;
  assign nS_st3_b237_c0 = nS_st2_b237_c0;
  assign nS_st3_b238_c0 = (nC_st2_b237_c0 == 0) ? nS_st2_b238_c0 : nS_st2_b238_c1;
  assign nS_st3_b239_c0 = (nC_st2_b237_c0 == 0) ? nS_st2_b239_c0 : nS_st2_b239_c1;
  assign nS_st3_b240_c0 = nS_st2_b240_c0;
  assign nS_st3_b241_c0 = nS_st2_b241_c0;
  assign nS_st3_b242_c0 = (nC_st2_b241_c0 == 0) ? nS_st2_b242_c0 : nS_st2_b242_c1;
  assign nS_st3_b243_c0 = (nC_st2_b241_c0 == 0) ? nS_st2_b243_c0 : nS_st2_b243_c1;
  assign nS_st3_b244_c0 = nS_st2_b244_c0;
  assign nS_st3_b245_c0 = nS_st2_b245_c0;
  assign nS_st3_b246_c0 = (nC_st2_b245_c0 == 0) ? nS_st2_b246_c0 : nS_st2_b246_c1;
  assign nS_st3_b247_c0 = (nC_st2_b245_c0 == 0) ? nS_st2_b247_c0 : nS_st2_b247_c1;
  assign nS_st3_b248_c0 = nS_st2_b248_c0;
  assign nS_st3_b249_c0 = nS_st2_b249_c0;
  assign nS_st3_b250_c0 = (nC_st2_b249_c0 == 0) ? nS_st2_b250_c0 : nS_st2_b250_c1;
  assign nS_st3_b251_c0 = (nC_st2_b249_c0 == 0) ? nS_st2_b251_c0 : nS_st2_b251_c1;
  assign nS_st3_b252_c0 = nS_st2_b252_c0;
  assign nS_st3_b253_c0 = nS_st2_b253_c0;
  assign nS_st3_b254_c0 = (nC_st2_b253_c0 == 0) ? nS_st2_b254_c0 : nS_st2_b254_c1;
  assign nS_st3_b255_c0 = (nC_st2_b253_c0 == 0) ? nS_st2_b255_c0 : nS_st2_b255_c1;
  assign nS_st3_b0_c1 = nS_st2_b0_c1;
  assign nS_st3_b1_c1 = nS_st2_b1_c1;
  assign nS_st3_b2_c1 = (nC_st2_b1_c1 == 0) ? nS_st2_b2_c0 : nS_st2_b2_c1;
  assign nS_st3_b3_c1 = (nC_st2_b1_c1 == 0) ? nS_st2_b3_c0 : nS_st2_b3_c1;
  assign nS_st3_b4_c1 = nS_st2_b4_c1;
  assign nS_st3_b5_c1 = nS_st2_b5_c1;
  assign nS_st3_b6_c1 = (nC_st2_b5_c1 == 0) ? nS_st2_b6_c0 : nS_st2_b6_c1;
  assign nS_st3_b7_c1 = (nC_st2_b5_c1 == 0) ? nS_st2_b7_c0 : nS_st2_b7_c1;
  assign nS_st3_b8_c1 = nS_st2_b8_c1;
  assign nS_st3_b9_c1 = nS_st2_b9_c1;
  assign nS_st3_b10_c1 = (nC_st2_b9_c1 == 0) ? nS_st2_b10_c0 : nS_st2_b10_c1;
  assign nS_st3_b11_c1 = (nC_st2_b9_c1 == 0) ? nS_st2_b11_c0 : nS_st2_b11_c1;
  assign nS_st3_b12_c1 = nS_st2_b12_c1;
  assign nS_st3_b13_c1 = nS_st2_b13_c1;
  assign nS_st3_b14_c1 = (nC_st2_b13_c1 == 0) ? nS_st2_b14_c0 : nS_st2_b14_c1;
  assign nS_st3_b15_c1 = (nC_st2_b13_c1 == 0) ? nS_st2_b15_c0 : nS_st2_b15_c1;
  assign nS_st3_b16_c1 = nS_st2_b16_c1;
  assign nS_st3_b17_c1 = nS_st2_b17_c1;
  assign nS_st3_b18_c1 = (nC_st2_b17_c1 == 0) ? nS_st2_b18_c0 : nS_st2_b18_c1;
  assign nS_st3_b19_c1 = (nC_st2_b17_c1 == 0) ? nS_st2_b19_c0 : nS_st2_b19_c1;
  assign nS_st3_b20_c1 = nS_st2_b20_c1;
  assign nS_st3_b21_c1 = nS_st2_b21_c1;
  assign nS_st3_b22_c1 = (nC_st2_b21_c1 == 0) ? nS_st2_b22_c0 : nS_st2_b22_c1;
  assign nS_st3_b23_c1 = (nC_st2_b21_c1 == 0) ? nS_st2_b23_c0 : nS_st2_b23_c1;
  assign nS_st3_b24_c1 = nS_st2_b24_c1;
  assign nS_st3_b25_c1 = nS_st2_b25_c1;
  assign nS_st3_b26_c1 = (nC_st2_b25_c1 == 0) ? nS_st2_b26_c0 : nS_st2_b26_c1;
  assign nS_st3_b27_c1 = (nC_st2_b25_c1 == 0) ? nS_st2_b27_c0 : nS_st2_b27_c1;
  assign nS_st3_b28_c1 = nS_st2_b28_c1;
  assign nS_st3_b29_c1 = nS_st2_b29_c1;
  assign nS_st3_b30_c1 = (nC_st2_b29_c1 == 0) ? nS_st2_b30_c0 : nS_st2_b30_c1;
  assign nS_st3_b31_c1 = (nC_st2_b29_c1 == 0) ? nS_st2_b31_c0 : nS_st2_b31_c1;
  assign nS_st3_b32_c1 = nS_st2_b32_c1;
  assign nS_st3_b33_c1 = nS_st2_b33_c1;
  assign nS_st3_b34_c1 = (nC_st2_b33_c1 == 0) ? nS_st2_b34_c0 : nS_st2_b34_c1;
  assign nS_st3_b35_c1 = (nC_st2_b33_c1 == 0) ? nS_st2_b35_c0 : nS_st2_b35_c1;
  assign nS_st3_b36_c1 = nS_st2_b36_c1;
  assign nS_st3_b37_c1 = nS_st2_b37_c1;
  assign nS_st3_b38_c1 = (nC_st2_b37_c1 == 0) ? nS_st2_b38_c0 : nS_st2_b38_c1;
  assign nS_st3_b39_c1 = (nC_st2_b37_c1 == 0) ? nS_st2_b39_c0 : nS_st2_b39_c1;
  assign nS_st3_b40_c1 = nS_st2_b40_c1;
  assign nS_st3_b41_c1 = nS_st2_b41_c1;
  assign nS_st3_b42_c1 = (nC_st2_b41_c1 == 0) ? nS_st2_b42_c0 : nS_st2_b42_c1;
  assign nS_st3_b43_c1 = (nC_st2_b41_c1 == 0) ? nS_st2_b43_c0 : nS_st2_b43_c1;
  assign nS_st3_b44_c1 = nS_st2_b44_c1;
  assign nS_st3_b45_c1 = nS_st2_b45_c1;
  assign nS_st3_b46_c1 = (nC_st2_b45_c1 == 0) ? nS_st2_b46_c0 : nS_st2_b46_c1;
  assign nS_st3_b47_c1 = (nC_st2_b45_c1 == 0) ? nS_st2_b47_c0 : nS_st2_b47_c1;
  assign nS_st3_b48_c1 = nS_st2_b48_c1;
  assign nS_st3_b49_c1 = nS_st2_b49_c1;
  assign nS_st3_b50_c1 = (nC_st2_b49_c1 == 0) ? nS_st2_b50_c0 : nS_st2_b50_c1;
  assign nS_st3_b51_c1 = (nC_st2_b49_c1 == 0) ? nS_st2_b51_c0 : nS_st2_b51_c1;
  assign nS_st3_b52_c1 = nS_st2_b52_c1;
  assign nS_st3_b53_c1 = nS_st2_b53_c1;
  assign nS_st3_b54_c1 = (nC_st2_b53_c1 == 0) ? nS_st2_b54_c0 : nS_st2_b54_c1;
  assign nS_st3_b55_c1 = (nC_st2_b53_c1 == 0) ? nS_st2_b55_c0 : nS_st2_b55_c1;
  assign nS_st3_b56_c1 = nS_st2_b56_c1;
  assign nS_st3_b57_c1 = nS_st2_b57_c1;
  assign nS_st3_b58_c1 = (nC_st2_b57_c1 == 0) ? nS_st2_b58_c0 : nS_st2_b58_c1;
  assign nS_st3_b59_c1 = (nC_st2_b57_c1 == 0) ? nS_st2_b59_c0 : nS_st2_b59_c1;
  assign nS_st3_b60_c1 = nS_st2_b60_c1;
  assign nS_st3_b61_c1 = nS_st2_b61_c1;
  assign nS_st3_b62_c1 = (nC_st2_b61_c1 == 0) ? nS_st2_b62_c0 : nS_st2_b62_c1;
  assign nS_st3_b63_c1 = (nC_st2_b61_c1 == 0) ? nS_st2_b63_c0 : nS_st2_b63_c1;
  assign nS_st3_b64_c1 = nS_st2_b64_c1;
  assign nS_st3_b65_c1 = nS_st2_b65_c1;
  assign nS_st3_b66_c1 = (nC_st2_b65_c1 == 0) ? nS_st2_b66_c0 : nS_st2_b66_c1;
  assign nS_st3_b67_c1 = (nC_st2_b65_c1 == 0) ? nS_st2_b67_c0 : nS_st2_b67_c1;
  assign nS_st3_b68_c1 = nS_st2_b68_c1;
  assign nS_st3_b69_c1 = nS_st2_b69_c1;
  assign nS_st3_b70_c1 = (nC_st2_b69_c1 == 0) ? nS_st2_b70_c0 : nS_st2_b70_c1;
  assign nS_st3_b71_c1 = (nC_st2_b69_c1 == 0) ? nS_st2_b71_c0 : nS_st2_b71_c1;
  assign nS_st3_b72_c1 = nS_st2_b72_c1;
  assign nS_st3_b73_c1 = nS_st2_b73_c1;
  assign nS_st3_b74_c1 = (nC_st2_b73_c1 == 0) ? nS_st2_b74_c0 : nS_st2_b74_c1;
  assign nS_st3_b75_c1 = (nC_st2_b73_c1 == 0) ? nS_st2_b75_c0 : nS_st2_b75_c1;
  assign nS_st3_b76_c1 = nS_st2_b76_c1;
  assign nS_st3_b77_c1 = nS_st2_b77_c1;
  assign nS_st3_b78_c1 = (nC_st2_b77_c1 == 0) ? nS_st2_b78_c0 : nS_st2_b78_c1;
  assign nS_st3_b79_c1 = (nC_st2_b77_c1 == 0) ? nS_st2_b79_c0 : nS_st2_b79_c1;
  assign nS_st3_b80_c1 = nS_st2_b80_c1;
  assign nS_st3_b81_c1 = nS_st2_b81_c1;
  assign nS_st3_b82_c1 = (nC_st2_b81_c1 == 0) ? nS_st2_b82_c0 : nS_st2_b82_c1;
  assign nS_st3_b83_c1 = (nC_st2_b81_c1 == 0) ? nS_st2_b83_c0 : nS_st2_b83_c1;
  assign nS_st3_b84_c1 = nS_st2_b84_c1;
  assign nS_st3_b85_c1 = nS_st2_b85_c1;
  assign nS_st3_b86_c1 = (nC_st2_b85_c1 == 0) ? nS_st2_b86_c0 : nS_st2_b86_c1;
  assign nS_st3_b87_c1 = (nC_st2_b85_c1 == 0) ? nS_st2_b87_c0 : nS_st2_b87_c1;
  assign nS_st3_b88_c1 = nS_st2_b88_c1;
  assign nS_st3_b89_c1 = nS_st2_b89_c1;
  assign nS_st3_b90_c1 = (nC_st2_b89_c1 == 0) ? nS_st2_b90_c0 : nS_st2_b90_c1;
  assign nS_st3_b91_c1 = (nC_st2_b89_c1 == 0) ? nS_st2_b91_c0 : nS_st2_b91_c1;
  assign nS_st3_b92_c1 = nS_st2_b92_c1;
  assign nS_st3_b93_c1 = nS_st2_b93_c1;
  assign nS_st3_b94_c1 = (nC_st2_b93_c1 == 0) ? nS_st2_b94_c0 : nS_st2_b94_c1;
  assign nS_st3_b95_c1 = (nC_st2_b93_c1 == 0) ? nS_st2_b95_c0 : nS_st2_b95_c1;
  assign nS_st3_b96_c1 = nS_st2_b96_c1;
  assign nS_st3_b97_c1 = nS_st2_b97_c1;
  assign nS_st3_b98_c1 = (nC_st2_b97_c1 == 0) ? nS_st2_b98_c0 : nS_st2_b98_c1;
  assign nS_st3_b99_c1 = (nC_st2_b97_c1 == 0) ? nS_st2_b99_c0 : nS_st2_b99_c1;
  assign nS_st3_b100_c1 = nS_st2_b100_c1;
  assign nS_st3_b101_c1 = nS_st2_b101_c1;
  assign nS_st3_b102_c1 = (nC_st2_b101_c1 == 0) ? nS_st2_b102_c0 : nS_st2_b102_c1;
  assign nS_st3_b103_c1 = (nC_st2_b101_c1 == 0) ? nS_st2_b103_c0 : nS_st2_b103_c1;
  assign nS_st3_b104_c1 = nS_st2_b104_c1;
  assign nS_st3_b105_c1 = nS_st2_b105_c1;
  assign nS_st3_b106_c1 = (nC_st2_b105_c1 == 0) ? nS_st2_b106_c0 : nS_st2_b106_c1;
  assign nS_st3_b107_c1 = (nC_st2_b105_c1 == 0) ? nS_st2_b107_c0 : nS_st2_b107_c1;
  assign nS_st3_b108_c1 = nS_st2_b108_c1;
  assign nS_st3_b109_c1 = nS_st2_b109_c1;
  assign nS_st3_b110_c1 = (nC_st2_b109_c1 == 0) ? nS_st2_b110_c0 : nS_st2_b110_c1;
  assign nS_st3_b111_c1 = (nC_st2_b109_c1 == 0) ? nS_st2_b111_c0 : nS_st2_b111_c1;
  assign nS_st3_b112_c1 = nS_st2_b112_c1;
  assign nS_st3_b113_c1 = nS_st2_b113_c1;
  assign nS_st3_b114_c1 = (nC_st2_b113_c1 == 0) ? nS_st2_b114_c0 : nS_st2_b114_c1;
  assign nS_st3_b115_c1 = (nC_st2_b113_c1 == 0) ? nS_st2_b115_c0 : nS_st2_b115_c1;
  assign nS_st3_b116_c1 = nS_st2_b116_c1;
  assign nS_st3_b117_c1 = nS_st2_b117_c1;
  assign nS_st3_b118_c1 = (nC_st2_b117_c1 == 0) ? nS_st2_b118_c0 : nS_st2_b118_c1;
  assign nS_st3_b119_c1 = (nC_st2_b117_c1 == 0) ? nS_st2_b119_c0 : nS_st2_b119_c1;
  assign nS_st3_b120_c1 = nS_st2_b120_c1;
  assign nS_st3_b121_c1 = nS_st2_b121_c1;
  assign nS_st3_b122_c1 = (nC_st2_b121_c1 == 0) ? nS_st2_b122_c0 : nS_st2_b122_c1;
  assign nS_st3_b123_c1 = (nC_st2_b121_c1 == 0) ? nS_st2_b123_c0 : nS_st2_b123_c1;
  assign nS_st3_b124_c1 = nS_st2_b124_c1;
  assign nS_st3_b125_c1 = nS_st2_b125_c1;
  assign nS_st3_b126_c1 = (nC_st2_b125_c1 == 0) ? nS_st2_b126_c0 : nS_st2_b126_c1;
  assign nS_st3_b127_c1 = (nC_st2_b125_c1 == 0) ? nS_st2_b127_c0 : nS_st2_b127_c1;
  assign nS_st3_b128_c1 = nS_st2_b128_c1;
  assign nS_st3_b129_c1 = nS_st2_b129_c1;
  assign nS_st3_b130_c1 = (nC_st2_b129_c1 == 0) ? nS_st2_b130_c0 : nS_st2_b130_c1;
  assign nS_st3_b131_c1 = (nC_st2_b129_c1 == 0) ? nS_st2_b131_c0 : nS_st2_b131_c1;
  assign nS_st3_b132_c1 = nS_st2_b132_c1;
  assign nS_st3_b133_c1 = nS_st2_b133_c1;
  assign nS_st3_b134_c1 = (nC_st2_b133_c1 == 0) ? nS_st2_b134_c0 : nS_st2_b134_c1;
  assign nS_st3_b135_c1 = (nC_st2_b133_c1 == 0) ? nS_st2_b135_c0 : nS_st2_b135_c1;
  assign nS_st3_b136_c1 = nS_st2_b136_c1;
  assign nS_st3_b137_c1 = nS_st2_b137_c1;
  assign nS_st3_b138_c1 = (nC_st2_b137_c1 == 0) ? nS_st2_b138_c0 : nS_st2_b138_c1;
  assign nS_st3_b139_c1 = (nC_st2_b137_c1 == 0) ? nS_st2_b139_c0 : nS_st2_b139_c1;
  assign nS_st3_b140_c1 = nS_st2_b140_c1;
  assign nS_st3_b141_c1 = nS_st2_b141_c1;
  assign nS_st3_b142_c1 = (nC_st2_b141_c1 == 0) ? nS_st2_b142_c0 : nS_st2_b142_c1;
  assign nS_st3_b143_c1 = (nC_st2_b141_c1 == 0) ? nS_st2_b143_c0 : nS_st2_b143_c1;
  assign nS_st3_b144_c1 = nS_st2_b144_c1;
  assign nS_st3_b145_c1 = nS_st2_b145_c1;
  assign nS_st3_b146_c1 = (nC_st2_b145_c1 == 0) ? nS_st2_b146_c0 : nS_st2_b146_c1;
  assign nS_st3_b147_c1 = (nC_st2_b145_c1 == 0) ? nS_st2_b147_c0 : nS_st2_b147_c1;
  assign nS_st3_b148_c1 = nS_st2_b148_c1;
  assign nS_st3_b149_c1 = nS_st2_b149_c1;
  assign nS_st3_b150_c1 = (nC_st2_b149_c1 == 0) ? nS_st2_b150_c0 : nS_st2_b150_c1;
  assign nS_st3_b151_c1 = (nC_st2_b149_c1 == 0) ? nS_st2_b151_c0 : nS_st2_b151_c1;
  assign nS_st3_b152_c1 = nS_st2_b152_c1;
  assign nS_st3_b153_c1 = nS_st2_b153_c1;
  assign nS_st3_b154_c1 = (nC_st2_b153_c1 == 0) ? nS_st2_b154_c0 : nS_st2_b154_c1;
  assign nS_st3_b155_c1 = (nC_st2_b153_c1 == 0) ? nS_st2_b155_c0 : nS_st2_b155_c1;
  assign nS_st3_b156_c1 = nS_st2_b156_c1;
  assign nS_st3_b157_c1 = nS_st2_b157_c1;
  assign nS_st3_b158_c1 = (nC_st2_b157_c1 == 0) ? nS_st2_b158_c0 : nS_st2_b158_c1;
  assign nS_st3_b159_c1 = (nC_st2_b157_c1 == 0) ? nS_st2_b159_c0 : nS_st2_b159_c1;
  assign nS_st3_b160_c1 = nS_st2_b160_c1;
  assign nS_st3_b161_c1 = nS_st2_b161_c1;
  assign nS_st3_b162_c1 = (nC_st2_b161_c1 == 0) ? nS_st2_b162_c0 : nS_st2_b162_c1;
  assign nS_st3_b163_c1 = (nC_st2_b161_c1 == 0) ? nS_st2_b163_c0 : nS_st2_b163_c1;
  assign nS_st3_b164_c1 = nS_st2_b164_c1;
  assign nS_st3_b165_c1 = nS_st2_b165_c1;
  assign nS_st3_b166_c1 = (nC_st2_b165_c1 == 0) ? nS_st2_b166_c0 : nS_st2_b166_c1;
  assign nS_st3_b167_c1 = (nC_st2_b165_c1 == 0) ? nS_st2_b167_c0 : nS_st2_b167_c1;
  assign nS_st3_b168_c1 = nS_st2_b168_c1;
  assign nS_st3_b169_c1 = nS_st2_b169_c1;
  assign nS_st3_b170_c1 = (nC_st2_b169_c1 == 0) ? nS_st2_b170_c0 : nS_st2_b170_c1;
  assign nS_st3_b171_c1 = (nC_st2_b169_c1 == 0) ? nS_st2_b171_c0 : nS_st2_b171_c1;
  assign nS_st3_b172_c1 = nS_st2_b172_c1;
  assign nS_st3_b173_c1 = nS_st2_b173_c1;
  assign nS_st3_b174_c1 = (nC_st2_b173_c1 == 0) ? nS_st2_b174_c0 : nS_st2_b174_c1;
  assign nS_st3_b175_c1 = (nC_st2_b173_c1 == 0) ? nS_st2_b175_c0 : nS_st2_b175_c1;
  assign nS_st3_b176_c1 = nS_st2_b176_c1;
  assign nS_st3_b177_c1 = nS_st2_b177_c1;
  assign nS_st3_b178_c1 = (nC_st2_b177_c1 == 0) ? nS_st2_b178_c0 : nS_st2_b178_c1;
  assign nS_st3_b179_c1 = (nC_st2_b177_c1 == 0) ? nS_st2_b179_c0 : nS_st2_b179_c1;
  assign nS_st3_b180_c1 = nS_st2_b180_c1;
  assign nS_st3_b181_c1 = nS_st2_b181_c1;
  assign nS_st3_b182_c1 = (nC_st2_b181_c1 == 0) ? nS_st2_b182_c0 : nS_st2_b182_c1;
  assign nS_st3_b183_c1 = (nC_st2_b181_c1 == 0) ? nS_st2_b183_c0 : nS_st2_b183_c1;
  assign nS_st3_b184_c1 = nS_st2_b184_c1;
  assign nS_st3_b185_c1 = nS_st2_b185_c1;
  assign nS_st3_b186_c1 = (nC_st2_b185_c1 == 0) ? nS_st2_b186_c0 : nS_st2_b186_c1;
  assign nS_st3_b187_c1 = (nC_st2_b185_c1 == 0) ? nS_st2_b187_c0 : nS_st2_b187_c1;
  assign nS_st3_b188_c1 = nS_st2_b188_c1;
  assign nS_st3_b189_c1 = nS_st2_b189_c1;
  assign nS_st3_b190_c1 = (nC_st2_b189_c1 == 0) ? nS_st2_b190_c0 : nS_st2_b190_c1;
  assign nS_st3_b191_c1 = (nC_st2_b189_c1 == 0) ? nS_st2_b191_c0 : nS_st2_b191_c1;
  assign nS_st3_b192_c1 = nS_st2_b192_c1;
  assign nS_st3_b193_c1 = nS_st2_b193_c1;
  assign nS_st3_b194_c1 = (nC_st2_b193_c1 == 0) ? nS_st2_b194_c0 : nS_st2_b194_c1;
  assign nS_st3_b195_c1 = (nC_st2_b193_c1 == 0) ? nS_st2_b195_c0 : nS_st2_b195_c1;
  assign nS_st3_b196_c1 = nS_st2_b196_c1;
  assign nS_st3_b197_c1 = nS_st2_b197_c1;
  assign nS_st3_b198_c1 = (nC_st2_b197_c1 == 0) ? nS_st2_b198_c0 : nS_st2_b198_c1;
  assign nS_st3_b199_c1 = (nC_st2_b197_c1 == 0) ? nS_st2_b199_c0 : nS_st2_b199_c1;
  assign nS_st3_b200_c1 = nS_st2_b200_c1;
  assign nS_st3_b201_c1 = nS_st2_b201_c1;
  assign nS_st3_b202_c1 = (nC_st2_b201_c1 == 0) ? nS_st2_b202_c0 : nS_st2_b202_c1;
  assign nS_st3_b203_c1 = (nC_st2_b201_c1 == 0) ? nS_st2_b203_c0 : nS_st2_b203_c1;
  assign nS_st3_b204_c1 = nS_st2_b204_c1;
  assign nS_st3_b205_c1 = nS_st2_b205_c1;
  assign nS_st3_b206_c1 = (nC_st2_b205_c1 == 0) ? nS_st2_b206_c0 : nS_st2_b206_c1;
  assign nS_st3_b207_c1 = (nC_st2_b205_c1 == 0) ? nS_st2_b207_c0 : nS_st2_b207_c1;
  assign nS_st3_b208_c1 = nS_st2_b208_c1;
  assign nS_st3_b209_c1 = nS_st2_b209_c1;
  assign nS_st3_b210_c1 = (nC_st2_b209_c1 == 0) ? nS_st2_b210_c0 : nS_st2_b210_c1;
  assign nS_st3_b211_c1 = (nC_st2_b209_c1 == 0) ? nS_st2_b211_c0 : nS_st2_b211_c1;
  assign nS_st3_b212_c1 = nS_st2_b212_c1;
  assign nS_st3_b213_c1 = nS_st2_b213_c1;
  assign nS_st3_b214_c1 = (nC_st2_b213_c1 == 0) ? nS_st2_b214_c0 : nS_st2_b214_c1;
  assign nS_st3_b215_c1 = (nC_st2_b213_c1 == 0) ? nS_st2_b215_c0 : nS_st2_b215_c1;
  assign nS_st3_b216_c1 = nS_st2_b216_c1;
  assign nS_st3_b217_c1 = nS_st2_b217_c1;
  assign nS_st3_b218_c1 = (nC_st2_b217_c1 == 0) ? nS_st2_b218_c0 : nS_st2_b218_c1;
  assign nS_st3_b219_c1 = (nC_st2_b217_c1 == 0) ? nS_st2_b219_c0 : nS_st2_b219_c1;
  assign nS_st3_b220_c1 = nS_st2_b220_c1;
  assign nS_st3_b221_c1 = nS_st2_b221_c1;
  assign nS_st3_b222_c1 = (nC_st2_b221_c1 == 0) ? nS_st2_b222_c0 : nS_st2_b222_c1;
  assign nS_st3_b223_c1 = (nC_st2_b221_c1 == 0) ? nS_st2_b223_c0 : nS_st2_b223_c1;
  assign nS_st3_b224_c1 = nS_st2_b224_c1;
  assign nS_st3_b225_c1 = nS_st2_b225_c1;
  assign nS_st3_b226_c1 = (nC_st2_b225_c1 == 0) ? nS_st2_b226_c0 : nS_st2_b226_c1;
  assign nS_st3_b227_c1 = (nC_st2_b225_c1 == 0) ? nS_st2_b227_c0 : nS_st2_b227_c1;
  assign nS_st3_b228_c1 = nS_st2_b228_c1;
  assign nS_st3_b229_c1 = nS_st2_b229_c1;
  assign nS_st3_b230_c1 = (nC_st2_b229_c1 == 0) ? nS_st2_b230_c0 : nS_st2_b230_c1;
  assign nS_st3_b231_c1 = (nC_st2_b229_c1 == 0) ? nS_st2_b231_c0 : nS_st2_b231_c1;
  assign nS_st3_b232_c1 = nS_st2_b232_c1;
  assign nS_st3_b233_c1 = nS_st2_b233_c1;
  assign nS_st3_b234_c1 = (nC_st2_b233_c1 == 0) ? nS_st2_b234_c0 : nS_st2_b234_c1;
  assign nS_st3_b235_c1 = (nC_st2_b233_c1 == 0) ? nS_st2_b235_c0 : nS_st2_b235_c1;
  assign nS_st3_b236_c1 = nS_st2_b236_c1;
  assign nS_st3_b237_c1 = nS_st2_b237_c1;
  assign nS_st3_b238_c1 = (nC_st2_b237_c1 == 0) ? nS_st2_b238_c0 : nS_st2_b238_c1;
  assign nS_st3_b239_c1 = (nC_st2_b237_c1 == 0) ? nS_st2_b239_c0 : nS_st2_b239_c1;
  assign nS_st3_b240_c1 = nS_st2_b240_c1;
  assign nS_st3_b241_c1 = nS_st2_b241_c1;
  assign nS_st3_b242_c1 = (nC_st2_b241_c1 == 0) ? nS_st2_b242_c0 : nS_st2_b242_c1;
  assign nS_st3_b243_c1 = (nC_st2_b241_c1 == 0) ? nS_st2_b243_c0 : nS_st2_b243_c1;
  assign nS_st3_b244_c1 = nS_st2_b244_c1;
  assign nS_st3_b245_c1 = nS_st2_b245_c1;
  assign nS_st3_b246_c1 = (nC_st2_b245_c1 == 0) ? nS_st2_b246_c0 : nS_st2_b246_c1;
  assign nS_st3_b247_c1 = (nC_st2_b245_c1 == 0) ? nS_st2_b247_c0 : nS_st2_b247_c1;
  assign nS_st3_b248_c1 = nS_st2_b248_c1;
  assign nS_st3_b249_c1 = nS_st2_b249_c1;
  assign nS_st3_b250_c1 = (nC_st2_b249_c1 == 0) ? nS_st2_b250_c0 : nS_st2_b250_c1;
  assign nS_st3_b251_c1 = (nC_st2_b249_c1 == 0) ? nS_st2_b251_c0 : nS_st2_b251_c1;
  assign nS_st3_b252_c1 = nS_st2_b252_c1;
  assign nS_st3_b253_c1 = nS_st2_b253_c1;
  assign nS_st3_b254_c1 = (nC_st2_b253_c1 == 0) ? nS_st2_b254_c0 : nS_st2_b254_c1;
  assign nS_st3_b255_c1 = (nC_st2_b253_c1 == 0) ? nS_st2_b255_c0 : nS_st2_b255_c1;
  assign nC_st3_b3_c0 = (nC_st2_b1_c0 == 0) ? nC_st2_b3_c0 : nC_st2_b3_c1;
  assign nC_st3_b7_c0 = (nC_st2_b5_c0 == 0) ? nC_st2_b7_c0 : nC_st2_b7_c1;
  assign nC_st3_b11_c0 = (nC_st2_b9_c0 == 0) ? nC_st2_b11_c0 : nC_st2_b11_c1;
  assign nC_st3_b15_c0 = (nC_st2_b13_c0 == 0) ? nC_st2_b15_c0 : nC_st2_b15_c1;
  assign nC_st3_b19_c0 = (nC_st2_b17_c0 == 0) ? nC_st2_b19_c0 : nC_st2_b19_c1;
  assign nC_st3_b23_c0 = (nC_st2_b21_c0 == 0) ? nC_st2_b23_c0 : nC_st2_b23_c1;
  assign nC_st3_b27_c0 = (nC_st2_b25_c0 == 0) ? nC_st2_b27_c0 : nC_st2_b27_c1;
  assign nC_st3_b31_c0 = (nC_st2_b29_c0 == 0) ? nC_st2_b31_c0 : nC_st2_b31_c1;
  assign nC_st3_b35_c0 = (nC_st2_b33_c0 == 0) ? nC_st2_b35_c0 : nC_st2_b35_c1;
  assign nC_st3_b39_c0 = (nC_st2_b37_c0 == 0) ? nC_st2_b39_c0 : nC_st2_b39_c1;
  assign nC_st3_b43_c0 = (nC_st2_b41_c0 == 0) ? nC_st2_b43_c0 : nC_st2_b43_c1;
  assign nC_st3_b47_c0 = (nC_st2_b45_c0 == 0) ? nC_st2_b47_c0 : nC_st2_b47_c1;
  assign nC_st3_b51_c0 = (nC_st2_b49_c0 == 0) ? nC_st2_b51_c0 : nC_st2_b51_c1;
  assign nC_st3_b55_c0 = (nC_st2_b53_c0 == 0) ? nC_st2_b55_c0 : nC_st2_b55_c1;
  assign nC_st3_b59_c0 = (nC_st2_b57_c0 == 0) ? nC_st2_b59_c0 : nC_st2_b59_c1;
  assign nC_st3_b63_c0 = (nC_st2_b61_c0 == 0) ? nC_st2_b63_c0 : nC_st2_b63_c1;
  assign nC_st3_b67_c0 = (nC_st2_b65_c0 == 0) ? nC_st2_b67_c0 : nC_st2_b67_c1;
  assign nC_st3_b71_c0 = (nC_st2_b69_c0 == 0) ? nC_st2_b71_c0 : nC_st2_b71_c1;
  assign nC_st3_b75_c0 = (nC_st2_b73_c0 == 0) ? nC_st2_b75_c0 : nC_st2_b75_c1;
  assign nC_st3_b79_c0 = (nC_st2_b77_c0 == 0) ? nC_st2_b79_c0 : nC_st2_b79_c1;
  assign nC_st3_b83_c0 = (nC_st2_b81_c0 == 0) ? nC_st2_b83_c0 : nC_st2_b83_c1;
  assign nC_st3_b87_c0 = (nC_st2_b85_c0 == 0) ? nC_st2_b87_c0 : nC_st2_b87_c1;
  assign nC_st3_b91_c0 = (nC_st2_b89_c0 == 0) ? nC_st2_b91_c0 : nC_st2_b91_c1;
  assign nC_st3_b95_c0 = (nC_st2_b93_c0 == 0) ? nC_st2_b95_c0 : nC_st2_b95_c1;
  assign nC_st3_b99_c0 = (nC_st2_b97_c0 == 0) ? nC_st2_b99_c0 : nC_st2_b99_c1;
  assign nC_st3_b103_c0 = (nC_st2_b101_c0 == 0) ? nC_st2_b103_c0 : nC_st2_b103_c1;
  assign nC_st3_b107_c0 = (nC_st2_b105_c0 == 0) ? nC_st2_b107_c0 : nC_st2_b107_c1;
  assign nC_st3_b111_c0 = (nC_st2_b109_c0 == 0) ? nC_st2_b111_c0 : nC_st2_b111_c1;
  assign nC_st3_b115_c0 = (nC_st2_b113_c0 == 0) ? nC_st2_b115_c0 : nC_st2_b115_c1;
  assign nC_st3_b119_c0 = (nC_st2_b117_c0 == 0) ? nC_st2_b119_c0 : nC_st2_b119_c1;
  assign nC_st3_b123_c0 = (nC_st2_b121_c0 == 0) ? nC_st2_b123_c0 : nC_st2_b123_c1;
  assign nC_st3_b127_c0 = (nC_st2_b125_c0 == 0) ? nC_st2_b127_c0 : nC_st2_b127_c1;
  assign nC_st3_b131_c0 = (nC_st2_b129_c0 == 0) ? nC_st2_b131_c0 : nC_st2_b131_c1;
  assign nC_st3_b135_c0 = (nC_st2_b133_c0 == 0) ? nC_st2_b135_c0 : nC_st2_b135_c1;
  assign nC_st3_b139_c0 = (nC_st2_b137_c0 == 0) ? nC_st2_b139_c0 : nC_st2_b139_c1;
  assign nC_st3_b143_c0 = (nC_st2_b141_c0 == 0) ? nC_st2_b143_c0 : nC_st2_b143_c1;
  assign nC_st3_b147_c0 = (nC_st2_b145_c0 == 0) ? nC_st2_b147_c0 : nC_st2_b147_c1;
  assign nC_st3_b151_c0 = (nC_st2_b149_c0 == 0) ? nC_st2_b151_c0 : nC_st2_b151_c1;
  assign nC_st3_b155_c0 = (nC_st2_b153_c0 == 0) ? nC_st2_b155_c0 : nC_st2_b155_c1;
  assign nC_st3_b159_c0 = (nC_st2_b157_c0 == 0) ? nC_st2_b159_c0 : nC_st2_b159_c1;
  assign nC_st3_b163_c0 = (nC_st2_b161_c0 == 0) ? nC_st2_b163_c0 : nC_st2_b163_c1;
  assign nC_st3_b167_c0 = (nC_st2_b165_c0 == 0) ? nC_st2_b167_c0 : nC_st2_b167_c1;
  assign nC_st3_b171_c0 = (nC_st2_b169_c0 == 0) ? nC_st2_b171_c0 : nC_st2_b171_c1;
  assign nC_st3_b175_c0 = (nC_st2_b173_c0 == 0) ? nC_st2_b175_c0 : nC_st2_b175_c1;
  assign nC_st3_b179_c0 = (nC_st2_b177_c0 == 0) ? nC_st2_b179_c0 : nC_st2_b179_c1;
  assign nC_st3_b183_c0 = (nC_st2_b181_c0 == 0) ? nC_st2_b183_c0 : nC_st2_b183_c1;
  assign nC_st3_b187_c0 = (nC_st2_b185_c0 == 0) ? nC_st2_b187_c0 : nC_st2_b187_c1;
  assign nC_st3_b191_c0 = (nC_st2_b189_c0 == 0) ? nC_st2_b191_c0 : nC_st2_b191_c1;
  assign nC_st3_b195_c0 = (nC_st2_b193_c0 == 0) ? nC_st2_b195_c0 : nC_st2_b195_c1;
  assign nC_st3_b199_c0 = (nC_st2_b197_c0 == 0) ? nC_st2_b199_c0 : nC_st2_b199_c1;
  assign nC_st3_b203_c0 = (nC_st2_b201_c0 == 0) ? nC_st2_b203_c0 : nC_st2_b203_c1;
  assign nC_st3_b207_c0 = (nC_st2_b205_c0 == 0) ? nC_st2_b207_c0 : nC_st2_b207_c1;
  assign nC_st3_b211_c0 = (nC_st2_b209_c0 == 0) ? nC_st2_b211_c0 : nC_st2_b211_c1;
  assign nC_st3_b215_c0 = (nC_st2_b213_c0 == 0) ? nC_st2_b215_c0 : nC_st2_b215_c1;
  assign nC_st3_b219_c0 = (nC_st2_b217_c0 == 0) ? nC_st2_b219_c0 : nC_st2_b219_c1;
  assign nC_st3_b223_c0 = (nC_st2_b221_c0 == 0) ? nC_st2_b223_c0 : nC_st2_b223_c1;
  assign nC_st3_b227_c0 = (nC_st2_b225_c0 == 0) ? nC_st2_b227_c0 : nC_st2_b227_c1;
  assign nC_st3_b231_c0 = (nC_st2_b229_c0 == 0) ? nC_st2_b231_c0 : nC_st2_b231_c1;
  assign nC_st3_b235_c0 = (nC_st2_b233_c0 == 0) ? nC_st2_b235_c0 : nC_st2_b235_c1;
  assign nC_st3_b239_c0 = (nC_st2_b237_c0 == 0) ? nC_st2_b239_c0 : nC_st2_b239_c1;
  assign nC_st3_b243_c0 = (nC_st2_b241_c0 == 0) ? nC_st2_b243_c0 : nC_st2_b243_c1;
  assign nC_st3_b247_c0 = (nC_st2_b245_c0 == 0) ? nC_st2_b247_c0 : nC_st2_b247_c1;
  assign nC_st3_b251_c0 = (nC_st2_b249_c0 == 0) ? nC_st2_b251_c0 : nC_st2_b251_c1;
  assign nC_st3_b255_c0 = (nC_st2_b253_c0 == 0) ? nC_st2_b255_c0 : nC_st2_b255_c1;
  assign nC_st3_b3_c1 = (nC_st2_b1_c1 == 0) ? nC_st2_b3_c0 : nC_st2_b3_c1;
  assign nC_st3_b7_c1 = (nC_st2_b5_c1 == 0) ? nC_st2_b7_c0 : nC_st2_b7_c1;
  assign nC_st3_b11_c1 = (nC_st2_b9_c1 == 0) ? nC_st2_b11_c0 : nC_st2_b11_c1;
  assign nC_st3_b15_c1 = (nC_st2_b13_c1 == 0) ? nC_st2_b15_c0 : nC_st2_b15_c1;
  assign nC_st3_b19_c1 = (nC_st2_b17_c1 == 0) ? nC_st2_b19_c0 : nC_st2_b19_c1;
  assign nC_st3_b23_c1 = (nC_st2_b21_c1 == 0) ? nC_st2_b23_c0 : nC_st2_b23_c1;
  assign nC_st3_b27_c1 = (nC_st2_b25_c1 == 0) ? nC_st2_b27_c0 : nC_st2_b27_c1;
  assign nC_st3_b31_c1 = (nC_st2_b29_c1 == 0) ? nC_st2_b31_c0 : nC_st2_b31_c1;
  assign nC_st3_b35_c1 = (nC_st2_b33_c1 == 0) ? nC_st2_b35_c0 : nC_st2_b35_c1;
  assign nC_st3_b39_c1 = (nC_st2_b37_c1 == 0) ? nC_st2_b39_c0 : nC_st2_b39_c1;
  assign nC_st3_b43_c1 = (nC_st2_b41_c1 == 0) ? nC_st2_b43_c0 : nC_st2_b43_c1;
  assign nC_st3_b47_c1 = (nC_st2_b45_c1 == 0) ? nC_st2_b47_c0 : nC_st2_b47_c1;
  assign nC_st3_b51_c1 = (nC_st2_b49_c1 == 0) ? nC_st2_b51_c0 : nC_st2_b51_c1;
  assign nC_st3_b55_c1 = (nC_st2_b53_c1 == 0) ? nC_st2_b55_c0 : nC_st2_b55_c1;
  assign nC_st3_b59_c1 = (nC_st2_b57_c1 == 0) ? nC_st2_b59_c0 : nC_st2_b59_c1;
  assign nC_st3_b63_c1 = (nC_st2_b61_c1 == 0) ? nC_st2_b63_c0 : nC_st2_b63_c1;
  assign nC_st3_b67_c1 = (nC_st2_b65_c1 == 0) ? nC_st2_b67_c0 : nC_st2_b67_c1;
  assign nC_st3_b71_c1 = (nC_st2_b69_c1 == 0) ? nC_st2_b71_c0 : nC_st2_b71_c1;
  assign nC_st3_b75_c1 = (nC_st2_b73_c1 == 0) ? nC_st2_b75_c0 : nC_st2_b75_c1;
  assign nC_st3_b79_c1 = (nC_st2_b77_c1 == 0) ? nC_st2_b79_c0 : nC_st2_b79_c1;
  assign nC_st3_b83_c1 = (nC_st2_b81_c1 == 0) ? nC_st2_b83_c0 : nC_st2_b83_c1;
  assign nC_st3_b87_c1 = (nC_st2_b85_c1 == 0) ? nC_st2_b87_c0 : nC_st2_b87_c1;
  assign nC_st3_b91_c1 = (nC_st2_b89_c1 == 0) ? nC_st2_b91_c0 : nC_st2_b91_c1;
  assign nC_st3_b95_c1 = (nC_st2_b93_c1 == 0) ? nC_st2_b95_c0 : nC_st2_b95_c1;
  assign nC_st3_b99_c1 = (nC_st2_b97_c1 == 0) ? nC_st2_b99_c0 : nC_st2_b99_c1;
  assign nC_st3_b103_c1 = (nC_st2_b101_c1 == 0) ? nC_st2_b103_c0 : nC_st2_b103_c1;
  assign nC_st3_b107_c1 = (nC_st2_b105_c1 == 0) ? nC_st2_b107_c0 : nC_st2_b107_c1;
  assign nC_st3_b111_c1 = (nC_st2_b109_c1 == 0) ? nC_st2_b111_c0 : nC_st2_b111_c1;
  assign nC_st3_b115_c1 = (nC_st2_b113_c1 == 0) ? nC_st2_b115_c0 : nC_st2_b115_c1;
  assign nC_st3_b119_c1 = (nC_st2_b117_c1 == 0) ? nC_st2_b119_c0 : nC_st2_b119_c1;
  assign nC_st3_b123_c1 = (nC_st2_b121_c1 == 0) ? nC_st2_b123_c0 : nC_st2_b123_c1;
  assign nC_st3_b127_c1 = (nC_st2_b125_c1 == 0) ? nC_st2_b127_c0 : nC_st2_b127_c1;
  assign nC_st3_b131_c1 = (nC_st2_b129_c1 == 0) ? nC_st2_b131_c0 : nC_st2_b131_c1;
  assign nC_st3_b135_c1 = (nC_st2_b133_c1 == 0) ? nC_st2_b135_c0 : nC_st2_b135_c1;
  assign nC_st3_b139_c1 = (nC_st2_b137_c1 == 0) ? nC_st2_b139_c0 : nC_st2_b139_c1;
  assign nC_st3_b143_c1 = (nC_st2_b141_c1 == 0) ? nC_st2_b143_c0 : nC_st2_b143_c1;
  assign nC_st3_b147_c1 = (nC_st2_b145_c1 == 0) ? nC_st2_b147_c0 : nC_st2_b147_c1;
  assign nC_st3_b151_c1 = (nC_st2_b149_c1 == 0) ? nC_st2_b151_c0 : nC_st2_b151_c1;
  assign nC_st3_b155_c1 = (nC_st2_b153_c1 == 0) ? nC_st2_b155_c0 : nC_st2_b155_c1;
  assign nC_st3_b159_c1 = (nC_st2_b157_c1 == 0) ? nC_st2_b159_c0 : nC_st2_b159_c1;
  assign nC_st3_b163_c1 = (nC_st2_b161_c1 == 0) ? nC_st2_b163_c0 : nC_st2_b163_c1;
  assign nC_st3_b167_c1 = (nC_st2_b165_c1 == 0) ? nC_st2_b167_c0 : nC_st2_b167_c1;
  assign nC_st3_b171_c1 = (nC_st2_b169_c1 == 0) ? nC_st2_b171_c0 : nC_st2_b171_c1;
  assign nC_st3_b175_c1 = (nC_st2_b173_c1 == 0) ? nC_st2_b175_c0 : nC_st2_b175_c1;
  assign nC_st3_b179_c1 = (nC_st2_b177_c1 == 0) ? nC_st2_b179_c0 : nC_st2_b179_c1;
  assign nC_st3_b183_c1 = (nC_st2_b181_c1 == 0) ? nC_st2_b183_c0 : nC_st2_b183_c1;
  assign nC_st3_b187_c1 = (nC_st2_b185_c1 == 0) ? nC_st2_b187_c0 : nC_st2_b187_c1;
  assign nC_st3_b191_c1 = (nC_st2_b189_c1 == 0) ? nC_st2_b191_c0 : nC_st2_b191_c1;
  assign nC_st3_b195_c1 = (nC_st2_b193_c1 == 0) ? nC_st2_b195_c0 : nC_st2_b195_c1;
  assign nC_st3_b199_c1 = (nC_st2_b197_c1 == 0) ? nC_st2_b199_c0 : nC_st2_b199_c1;
  assign nC_st3_b203_c1 = (nC_st2_b201_c1 == 0) ? nC_st2_b203_c0 : nC_st2_b203_c1;
  assign nC_st3_b207_c1 = (nC_st2_b205_c1 == 0) ? nC_st2_b207_c0 : nC_st2_b207_c1;
  assign nC_st3_b211_c1 = (nC_st2_b209_c1 == 0) ? nC_st2_b211_c0 : nC_st2_b211_c1;
  assign nC_st3_b215_c1 = (nC_st2_b213_c1 == 0) ? nC_st2_b215_c0 : nC_st2_b215_c1;
  assign nC_st3_b219_c1 = (nC_st2_b217_c1 == 0) ? nC_st2_b219_c0 : nC_st2_b219_c1;
  assign nC_st3_b223_c1 = (nC_st2_b221_c1 == 0) ? nC_st2_b223_c0 : nC_st2_b223_c1;
  assign nC_st3_b227_c1 = (nC_st2_b225_c1 == 0) ? nC_st2_b227_c0 : nC_st2_b227_c1;
  assign nC_st3_b231_c1 = (nC_st2_b229_c1 == 0) ? nC_st2_b231_c0 : nC_st2_b231_c1;
  assign nC_st3_b235_c1 = (nC_st2_b233_c1 == 0) ? nC_st2_b235_c0 : nC_st2_b235_c1;
  assign nC_st3_b239_c1 = (nC_st2_b237_c1 == 0) ? nC_st2_b239_c0 : nC_st2_b239_c1;
  assign nC_st3_b243_c1 = (nC_st2_b241_c1 == 0) ? nC_st2_b243_c0 : nC_st2_b243_c1;
  assign nC_st3_b247_c1 = (nC_st2_b245_c1 == 0) ? nC_st2_b247_c0 : nC_st2_b247_c1;
  assign nC_st3_b251_c1 = (nC_st2_b249_c1 == 0) ? nC_st2_b251_c0 : nC_st2_b251_c1;
  assign nC_st3_b255_c1 = (nC_st2_b253_c1 == 0) ? nC_st2_b255_c0 : nC_st2_b255_c1;

  assign nS_st4_b0_c0 = nS_st3_b0_c0;
  assign nS_st4_b1_c0 = nS_st3_b1_c0;
  assign nS_st4_b2_c0 = nS_st3_b2_c0;
  assign nS_st4_b3_c0 = nS_st3_b3_c0;
  assign nS_st4_b4_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b4_c0 : nS_st3_b4_c1;
  assign nS_st4_b5_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b5_c0 : nS_st3_b5_c1;
  assign nS_st4_b6_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b6_c0 : nS_st3_b6_c1;
  assign nS_st4_b7_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b7_c0 : nS_st3_b7_c1;
  assign nS_st4_b8_c0 = nS_st3_b8_c0;
  assign nS_st4_b9_c0 = nS_st3_b9_c0;
  assign nS_st4_b10_c0 = nS_st3_b10_c0;
  assign nS_st4_b11_c0 = nS_st3_b11_c0;
  assign nS_st4_b12_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b12_c0 : nS_st3_b12_c1;
  assign nS_st4_b13_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b13_c0 : nS_st3_b13_c1;
  assign nS_st4_b14_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b14_c0 : nS_st3_b14_c1;
  assign nS_st4_b15_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b15_c0 : nS_st3_b15_c1;
  assign nS_st4_b16_c0 = nS_st3_b16_c0;
  assign nS_st4_b17_c0 = nS_st3_b17_c0;
  assign nS_st4_b18_c0 = nS_st3_b18_c0;
  assign nS_st4_b19_c0 = nS_st3_b19_c0;
  assign nS_st4_b20_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b20_c0 : nS_st3_b20_c1;
  assign nS_st4_b21_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b21_c0 : nS_st3_b21_c1;
  assign nS_st4_b22_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b22_c0 : nS_st3_b22_c1;
  assign nS_st4_b23_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b23_c0 : nS_st3_b23_c1;
  assign nS_st4_b24_c0 = nS_st3_b24_c0;
  assign nS_st4_b25_c0 = nS_st3_b25_c0;
  assign nS_st4_b26_c0 = nS_st3_b26_c0;
  assign nS_st4_b27_c0 = nS_st3_b27_c0;
  assign nS_st4_b28_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b28_c0 : nS_st3_b28_c1;
  assign nS_st4_b29_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b29_c0 : nS_st3_b29_c1;
  assign nS_st4_b30_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b30_c0 : nS_st3_b30_c1;
  assign nS_st4_b31_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b31_c0 : nS_st3_b31_c1;
  assign nS_st4_b32_c0 = nS_st3_b32_c0;
  assign nS_st4_b33_c0 = nS_st3_b33_c0;
  assign nS_st4_b34_c0 = nS_st3_b34_c0;
  assign nS_st4_b35_c0 = nS_st3_b35_c0;
  assign nS_st4_b36_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b36_c0 : nS_st3_b36_c1;
  assign nS_st4_b37_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b37_c0 : nS_st3_b37_c1;
  assign nS_st4_b38_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b38_c0 : nS_st3_b38_c1;
  assign nS_st4_b39_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b39_c0 : nS_st3_b39_c1;
  assign nS_st4_b40_c0 = nS_st3_b40_c0;
  assign nS_st4_b41_c0 = nS_st3_b41_c0;
  assign nS_st4_b42_c0 = nS_st3_b42_c0;
  assign nS_st4_b43_c0 = nS_st3_b43_c0;
  assign nS_st4_b44_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b44_c0 : nS_st3_b44_c1;
  assign nS_st4_b45_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b45_c0 : nS_st3_b45_c1;
  assign nS_st4_b46_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b46_c0 : nS_st3_b46_c1;
  assign nS_st4_b47_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b47_c0 : nS_st3_b47_c1;
  assign nS_st4_b48_c0 = nS_st3_b48_c0;
  assign nS_st4_b49_c0 = nS_st3_b49_c0;
  assign nS_st4_b50_c0 = nS_st3_b50_c0;
  assign nS_st4_b51_c0 = nS_st3_b51_c0;
  assign nS_st4_b52_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b52_c0 : nS_st3_b52_c1;
  assign nS_st4_b53_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b53_c0 : nS_st3_b53_c1;
  assign nS_st4_b54_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b54_c0 : nS_st3_b54_c1;
  assign nS_st4_b55_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b55_c0 : nS_st3_b55_c1;
  assign nS_st4_b56_c0 = nS_st3_b56_c0;
  assign nS_st4_b57_c0 = nS_st3_b57_c0;
  assign nS_st4_b58_c0 = nS_st3_b58_c0;
  assign nS_st4_b59_c0 = nS_st3_b59_c0;
  assign nS_st4_b60_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b60_c0 : nS_st3_b60_c1;
  assign nS_st4_b61_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b61_c0 : nS_st3_b61_c1;
  assign nS_st4_b62_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b62_c0 : nS_st3_b62_c1;
  assign nS_st4_b63_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b63_c0 : nS_st3_b63_c1;
  assign nS_st4_b64_c0 = nS_st3_b64_c0;
  assign nS_st4_b65_c0 = nS_st3_b65_c0;
  assign nS_st4_b66_c0 = nS_st3_b66_c0;
  assign nS_st4_b67_c0 = nS_st3_b67_c0;
  assign nS_st4_b68_c0 = (nC_st3_b67_c0 == 0) ? nS_st3_b68_c0 : nS_st3_b68_c1;
  assign nS_st4_b69_c0 = (nC_st3_b67_c0 == 0) ? nS_st3_b69_c0 : nS_st3_b69_c1;
  assign nS_st4_b70_c0 = (nC_st3_b67_c0 == 0) ? nS_st3_b70_c0 : nS_st3_b70_c1;
  assign nS_st4_b71_c0 = (nC_st3_b67_c0 == 0) ? nS_st3_b71_c0 : nS_st3_b71_c1;
  assign nS_st4_b72_c0 = nS_st3_b72_c0;
  assign nS_st4_b73_c0 = nS_st3_b73_c0;
  assign nS_st4_b74_c0 = nS_st3_b74_c0;
  assign nS_st4_b75_c0 = nS_st3_b75_c0;
  assign nS_st4_b76_c0 = (nC_st3_b75_c0 == 0) ? nS_st3_b76_c0 : nS_st3_b76_c1;
  assign nS_st4_b77_c0 = (nC_st3_b75_c0 == 0) ? nS_st3_b77_c0 : nS_st3_b77_c1;
  assign nS_st4_b78_c0 = (nC_st3_b75_c0 == 0) ? nS_st3_b78_c0 : nS_st3_b78_c1;
  assign nS_st4_b79_c0 = (nC_st3_b75_c0 == 0) ? nS_st3_b79_c0 : nS_st3_b79_c1;
  assign nS_st4_b80_c0 = nS_st3_b80_c0;
  assign nS_st4_b81_c0 = nS_st3_b81_c0;
  assign nS_st4_b82_c0 = nS_st3_b82_c0;
  assign nS_st4_b83_c0 = nS_st3_b83_c0;
  assign nS_st4_b84_c0 = (nC_st3_b83_c0 == 0) ? nS_st3_b84_c0 : nS_st3_b84_c1;
  assign nS_st4_b85_c0 = (nC_st3_b83_c0 == 0) ? nS_st3_b85_c0 : nS_st3_b85_c1;
  assign nS_st4_b86_c0 = (nC_st3_b83_c0 == 0) ? nS_st3_b86_c0 : nS_st3_b86_c1;
  assign nS_st4_b87_c0 = (nC_st3_b83_c0 == 0) ? nS_st3_b87_c0 : nS_st3_b87_c1;
  assign nS_st4_b88_c0 = nS_st3_b88_c0;
  assign nS_st4_b89_c0 = nS_st3_b89_c0;
  assign nS_st4_b90_c0 = nS_st3_b90_c0;
  assign nS_st4_b91_c0 = nS_st3_b91_c0;
  assign nS_st4_b92_c0 = (nC_st3_b91_c0 == 0) ? nS_st3_b92_c0 : nS_st3_b92_c1;
  assign nS_st4_b93_c0 = (nC_st3_b91_c0 == 0) ? nS_st3_b93_c0 : nS_st3_b93_c1;
  assign nS_st4_b94_c0 = (nC_st3_b91_c0 == 0) ? nS_st3_b94_c0 : nS_st3_b94_c1;
  assign nS_st4_b95_c0 = (nC_st3_b91_c0 == 0) ? nS_st3_b95_c0 : nS_st3_b95_c1;
  assign nS_st4_b96_c0 = nS_st3_b96_c0;
  assign nS_st4_b97_c0 = nS_st3_b97_c0;
  assign nS_st4_b98_c0 = nS_st3_b98_c0;
  assign nS_st4_b99_c0 = nS_st3_b99_c0;
  assign nS_st4_b100_c0 = (nC_st3_b99_c0 == 0) ? nS_st3_b100_c0 : nS_st3_b100_c1;
  assign nS_st4_b101_c0 = (nC_st3_b99_c0 == 0) ? nS_st3_b101_c0 : nS_st3_b101_c1;
  assign nS_st4_b102_c0 = (nC_st3_b99_c0 == 0) ? nS_st3_b102_c0 : nS_st3_b102_c1;
  assign nS_st4_b103_c0 = (nC_st3_b99_c0 == 0) ? nS_st3_b103_c0 : nS_st3_b103_c1;
  assign nS_st4_b104_c0 = nS_st3_b104_c0;
  assign nS_st4_b105_c0 = nS_st3_b105_c0;
  assign nS_st4_b106_c0 = nS_st3_b106_c0;
  assign nS_st4_b107_c0 = nS_st3_b107_c0;
  assign nS_st4_b108_c0 = (nC_st3_b107_c0 == 0) ? nS_st3_b108_c0 : nS_st3_b108_c1;
  assign nS_st4_b109_c0 = (nC_st3_b107_c0 == 0) ? nS_st3_b109_c0 : nS_st3_b109_c1;
  assign nS_st4_b110_c0 = (nC_st3_b107_c0 == 0) ? nS_st3_b110_c0 : nS_st3_b110_c1;
  assign nS_st4_b111_c0 = (nC_st3_b107_c0 == 0) ? nS_st3_b111_c0 : nS_st3_b111_c1;
  assign nS_st4_b112_c0 = nS_st3_b112_c0;
  assign nS_st4_b113_c0 = nS_st3_b113_c0;
  assign nS_st4_b114_c0 = nS_st3_b114_c0;
  assign nS_st4_b115_c0 = nS_st3_b115_c0;
  assign nS_st4_b116_c0 = (nC_st3_b115_c0 == 0) ? nS_st3_b116_c0 : nS_st3_b116_c1;
  assign nS_st4_b117_c0 = (nC_st3_b115_c0 == 0) ? nS_st3_b117_c0 : nS_st3_b117_c1;
  assign nS_st4_b118_c0 = (nC_st3_b115_c0 == 0) ? nS_st3_b118_c0 : nS_st3_b118_c1;
  assign nS_st4_b119_c0 = (nC_st3_b115_c0 == 0) ? nS_st3_b119_c0 : nS_st3_b119_c1;
  assign nS_st4_b120_c0 = nS_st3_b120_c0;
  assign nS_st4_b121_c0 = nS_st3_b121_c0;
  assign nS_st4_b122_c0 = nS_st3_b122_c0;
  assign nS_st4_b123_c0 = nS_st3_b123_c0;
  assign nS_st4_b124_c0 = (nC_st3_b123_c0 == 0) ? nS_st3_b124_c0 : nS_st3_b124_c1;
  assign nS_st4_b125_c0 = (nC_st3_b123_c0 == 0) ? nS_st3_b125_c0 : nS_st3_b125_c1;
  assign nS_st4_b126_c0 = (nC_st3_b123_c0 == 0) ? nS_st3_b126_c0 : nS_st3_b126_c1;
  assign nS_st4_b127_c0 = (nC_st3_b123_c0 == 0) ? nS_st3_b127_c0 : nS_st3_b127_c1;
  assign nS_st4_b128_c0 = nS_st3_b128_c0;
  assign nS_st4_b129_c0 = nS_st3_b129_c0;
  assign nS_st4_b130_c0 = nS_st3_b130_c0;
  assign nS_st4_b131_c0 = nS_st3_b131_c0;
  assign nS_st4_b132_c0 = (nC_st3_b131_c0 == 0) ? nS_st3_b132_c0 : nS_st3_b132_c1;
  assign nS_st4_b133_c0 = (nC_st3_b131_c0 == 0) ? nS_st3_b133_c0 : nS_st3_b133_c1;
  assign nS_st4_b134_c0 = (nC_st3_b131_c0 == 0) ? nS_st3_b134_c0 : nS_st3_b134_c1;
  assign nS_st4_b135_c0 = (nC_st3_b131_c0 == 0) ? nS_st3_b135_c0 : nS_st3_b135_c1;
  assign nS_st4_b136_c0 = nS_st3_b136_c0;
  assign nS_st4_b137_c0 = nS_st3_b137_c0;
  assign nS_st4_b138_c0 = nS_st3_b138_c0;
  assign nS_st4_b139_c0 = nS_st3_b139_c0;
  assign nS_st4_b140_c0 = (nC_st3_b139_c0 == 0) ? nS_st3_b140_c0 : nS_st3_b140_c1;
  assign nS_st4_b141_c0 = (nC_st3_b139_c0 == 0) ? nS_st3_b141_c0 : nS_st3_b141_c1;
  assign nS_st4_b142_c0 = (nC_st3_b139_c0 == 0) ? nS_st3_b142_c0 : nS_st3_b142_c1;
  assign nS_st4_b143_c0 = (nC_st3_b139_c0 == 0) ? nS_st3_b143_c0 : nS_st3_b143_c1;
  assign nS_st4_b144_c0 = nS_st3_b144_c0;
  assign nS_st4_b145_c0 = nS_st3_b145_c0;
  assign nS_st4_b146_c0 = nS_st3_b146_c0;
  assign nS_st4_b147_c0 = nS_st3_b147_c0;
  assign nS_st4_b148_c0 = (nC_st3_b147_c0 == 0) ? nS_st3_b148_c0 : nS_st3_b148_c1;
  assign nS_st4_b149_c0 = (nC_st3_b147_c0 == 0) ? nS_st3_b149_c0 : nS_st3_b149_c1;
  assign nS_st4_b150_c0 = (nC_st3_b147_c0 == 0) ? nS_st3_b150_c0 : nS_st3_b150_c1;
  assign nS_st4_b151_c0 = (nC_st3_b147_c0 == 0) ? nS_st3_b151_c0 : nS_st3_b151_c1;
  assign nS_st4_b152_c0 = nS_st3_b152_c0;
  assign nS_st4_b153_c0 = nS_st3_b153_c0;
  assign nS_st4_b154_c0 = nS_st3_b154_c0;
  assign nS_st4_b155_c0 = nS_st3_b155_c0;
  assign nS_st4_b156_c0 = (nC_st3_b155_c0 == 0) ? nS_st3_b156_c0 : nS_st3_b156_c1;
  assign nS_st4_b157_c0 = (nC_st3_b155_c0 == 0) ? nS_st3_b157_c0 : nS_st3_b157_c1;
  assign nS_st4_b158_c0 = (nC_st3_b155_c0 == 0) ? nS_st3_b158_c0 : nS_st3_b158_c1;
  assign nS_st4_b159_c0 = (nC_st3_b155_c0 == 0) ? nS_st3_b159_c0 : nS_st3_b159_c1;
  assign nS_st4_b160_c0 = nS_st3_b160_c0;
  assign nS_st4_b161_c0 = nS_st3_b161_c0;
  assign nS_st4_b162_c0 = nS_st3_b162_c0;
  assign nS_st4_b163_c0 = nS_st3_b163_c0;
  assign nS_st4_b164_c0 = (nC_st3_b163_c0 == 0) ? nS_st3_b164_c0 : nS_st3_b164_c1;
  assign nS_st4_b165_c0 = (nC_st3_b163_c0 == 0) ? nS_st3_b165_c0 : nS_st3_b165_c1;
  assign nS_st4_b166_c0 = (nC_st3_b163_c0 == 0) ? nS_st3_b166_c0 : nS_st3_b166_c1;
  assign nS_st4_b167_c0 = (nC_st3_b163_c0 == 0) ? nS_st3_b167_c0 : nS_st3_b167_c1;
  assign nS_st4_b168_c0 = nS_st3_b168_c0;
  assign nS_st4_b169_c0 = nS_st3_b169_c0;
  assign nS_st4_b170_c0 = nS_st3_b170_c0;
  assign nS_st4_b171_c0 = nS_st3_b171_c0;
  assign nS_st4_b172_c0 = (nC_st3_b171_c0 == 0) ? nS_st3_b172_c0 : nS_st3_b172_c1;
  assign nS_st4_b173_c0 = (nC_st3_b171_c0 == 0) ? nS_st3_b173_c0 : nS_st3_b173_c1;
  assign nS_st4_b174_c0 = (nC_st3_b171_c0 == 0) ? nS_st3_b174_c0 : nS_st3_b174_c1;
  assign nS_st4_b175_c0 = (nC_st3_b171_c0 == 0) ? nS_st3_b175_c0 : nS_st3_b175_c1;
  assign nS_st4_b176_c0 = nS_st3_b176_c0;
  assign nS_st4_b177_c0 = nS_st3_b177_c0;
  assign nS_st4_b178_c0 = nS_st3_b178_c0;
  assign nS_st4_b179_c0 = nS_st3_b179_c0;
  assign nS_st4_b180_c0 = (nC_st3_b179_c0 == 0) ? nS_st3_b180_c0 : nS_st3_b180_c1;
  assign nS_st4_b181_c0 = (nC_st3_b179_c0 == 0) ? nS_st3_b181_c0 : nS_st3_b181_c1;
  assign nS_st4_b182_c0 = (nC_st3_b179_c0 == 0) ? nS_st3_b182_c0 : nS_st3_b182_c1;
  assign nS_st4_b183_c0 = (nC_st3_b179_c0 == 0) ? nS_st3_b183_c0 : nS_st3_b183_c1;
  assign nS_st4_b184_c0 = nS_st3_b184_c0;
  assign nS_st4_b185_c0 = nS_st3_b185_c0;
  assign nS_st4_b186_c0 = nS_st3_b186_c0;
  assign nS_st4_b187_c0 = nS_st3_b187_c0;
  assign nS_st4_b188_c0 = (nC_st3_b187_c0 == 0) ? nS_st3_b188_c0 : nS_st3_b188_c1;
  assign nS_st4_b189_c0 = (nC_st3_b187_c0 == 0) ? nS_st3_b189_c0 : nS_st3_b189_c1;
  assign nS_st4_b190_c0 = (nC_st3_b187_c0 == 0) ? nS_st3_b190_c0 : nS_st3_b190_c1;
  assign nS_st4_b191_c0 = (nC_st3_b187_c0 == 0) ? nS_st3_b191_c0 : nS_st3_b191_c1;
  assign nS_st4_b192_c0 = nS_st3_b192_c0;
  assign nS_st4_b193_c0 = nS_st3_b193_c0;
  assign nS_st4_b194_c0 = nS_st3_b194_c0;
  assign nS_st4_b195_c0 = nS_st3_b195_c0;
  assign nS_st4_b196_c0 = (nC_st3_b195_c0 == 0) ? nS_st3_b196_c0 : nS_st3_b196_c1;
  assign nS_st4_b197_c0 = (nC_st3_b195_c0 == 0) ? nS_st3_b197_c0 : nS_st3_b197_c1;
  assign nS_st4_b198_c0 = (nC_st3_b195_c0 == 0) ? nS_st3_b198_c0 : nS_st3_b198_c1;
  assign nS_st4_b199_c0 = (nC_st3_b195_c0 == 0) ? nS_st3_b199_c0 : nS_st3_b199_c1;
  assign nS_st4_b200_c0 = nS_st3_b200_c0;
  assign nS_st4_b201_c0 = nS_st3_b201_c0;
  assign nS_st4_b202_c0 = nS_st3_b202_c0;
  assign nS_st4_b203_c0 = nS_st3_b203_c0;
  assign nS_st4_b204_c0 = (nC_st3_b203_c0 == 0) ? nS_st3_b204_c0 : nS_st3_b204_c1;
  assign nS_st4_b205_c0 = (nC_st3_b203_c0 == 0) ? nS_st3_b205_c0 : nS_st3_b205_c1;
  assign nS_st4_b206_c0 = (nC_st3_b203_c0 == 0) ? nS_st3_b206_c0 : nS_st3_b206_c1;
  assign nS_st4_b207_c0 = (nC_st3_b203_c0 == 0) ? nS_st3_b207_c0 : nS_st3_b207_c1;
  assign nS_st4_b208_c0 = nS_st3_b208_c0;
  assign nS_st4_b209_c0 = nS_st3_b209_c0;
  assign nS_st4_b210_c0 = nS_st3_b210_c0;
  assign nS_st4_b211_c0 = nS_st3_b211_c0;
  assign nS_st4_b212_c0 = (nC_st3_b211_c0 == 0) ? nS_st3_b212_c0 : nS_st3_b212_c1;
  assign nS_st4_b213_c0 = (nC_st3_b211_c0 == 0) ? nS_st3_b213_c0 : nS_st3_b213_c1;
  assign nS_st4_b214_c0 = (nC_st3_b211_c0 == 0) ? nS_st3_b214_c0 : nS_st3_b214_c1;
  assign nS_st4_b215_c0 = (nC_st3_b211_c0 == 0) ? nS_st3_b215_c0 : nS_st3_b215_c1;
  assign nS_st4_b216_c0 = nS_st3_b216_c0;
  assign nS_st4_b217_c0 = nS_st3_b217_c0;
  assign nS_st4_b218_c0 = nS_st3_b218_c0;
  assign nS_st4_b219_c0 = nS_st3_b219_c0;
  assign nS_st4_b220_c0 = (nC_st3_b219_c0 == 0) ? nS_st3_b220_c0 : nS_st3_b220_c1;
  assign nS_st4_b221_c0 = (nC_st3_b219_c0 == 0) ? nS_st3_b221_c0 : nS_st3_b221_c1;
  assign nS_st4_b222_c0 = (nC_st3_b219_c0 == 0) ? nS_st3_b222_c0 : nS_st3_b222_c1;
  assign nS_st4_b223_c0 = (nC_st3_b219_c0 == 0) ? nS_st3_b223_c0 : nS_st3_b223_c1;
  assign nS_st4_b224_c0 = nS_st3_b224_c0;
  assign nS_st4_b225_c0 = nS_st3_b225_c0;
  assign nS_st4_b226_c0 = nS_st3_b226_c0;
  assign nS_st4_b227_c0 = nS_st3_b227_c0;
  assign nS_st4_b228_c0 = (nC_st3_b227_c0 == 0) ? nS_st3_b228_c0 : nS_st3_b228_c1;
  assign nS_st4_b229_c0 = (nC_st3_b227_c0 == 0) ? nS_st3_b229_c0 : nS_st3_b229_c1;
  assign nS_st4_b230_c0 = (nC_st3_b227_c0 == 0) ? nS_st3_b230_c0 : nS_st3_b230_c1;
  assign nS_st4_b231_c0 = (nC_st3_b227_c0 == 0) ? nS_st3_b231_c0 : nS_st3_b231_c1;
  assign nS_st4_b232_c0 = nS_st3_b232_c0;
  assign nS_st4_b233_c0 = nS_st3_b233_c0;
  assign nS_st4_b234_c0 = nS_st3_b234_c0;
  assign nS_st4_b235_c0 = nS_st3_b235_c0;
  assign nS_st4_b236_c0 = (nC_st3_b235_c0 == 0) ? nS_st3_b236_c0 : nS_st3_b236_c1;
  assign nS_st4_b237_c0 = (nC_st3_b235_c0 == 0) ? nS_st3_b237_c0 : nS_st3_b237_c1;
  assign nS_st4_b238_c0 = (nC_st3_b235_c0 == 0) ? nS_st3_b238_c0 : nS_st3_b238_c1;
  assign nS_st4_b239_c0 = (nC_st3_b235_c0 == 0) ? nS_st3_b239_c0 : nS_st3_b239_c1;
  assign nS_st4_b240_c0 = nS_st3_b240_c0;
  assign nS_st4_b241_c0 = nS_st3_b241_c0;
  assign nS_st4_b242_c0 = nS_st3_b242_c0;
  assign nS_st4_b243_c0 = nS_st3_b243_c0;
  assign nS_st4_b244_c0 = (nC_st3_b243_c0 == 0) ? nS_st3_b244_c0 : nS_st3_b244_c1;
  assign nS_st4_b245_c0 = (nC_st3_b243_c0 == 0) ? nS_st3_b245_c0 : nS_st3_b245_c1;
  assign nS_st4_b246_c0 = (nC_st3_b243_c0 == 0) ? nS_st3_b246_c0 : nS_st3_b246_c1;
  assign nS_st4_b247_c0 = (nC_st3_b243_c0 == 0) ? nS_st3_b247_c0 : nS_st3_b247_c1;
  assign nS_st4_b248_c0 = nS_st3_b248_c0;
  assign nS_st4_b249_c0 = nS_st3_b249_c0;
  assign nS_st4_b250_c0 = nS_st3_b250_c0;
  assign nS_st4_b251_c0 = nS_st3_b251_c0;
  assign nS_st4_b252_c0 = (nC_st3_b251_c0 == 0) ? nS_st3_b252_c0 : nS_st3_b252_c1;
  assign nS_st4_b253_c0 = (nC_st3_b251_c0 == 0) ? nS_st3_b253_c0 : nS_st3_b253_c1;
  assign nS_st4_b254_c0 = (nC_st3_b251_c0 == 0) ? nS_st3_b254_c0 : nS_st3_b254_c1;
  assign nS_st4_b255_c0 = (nC_st3_b251_c0 == 0) ? nS_st3_b255_c0 : nS_st3_b255_c1;
  assign nS_st4_b0_c1 = nS_st3_b0_c1;
  assign nS_st4_b1_c1 = nS_st3_b1_c1;
  assign nS_st4_b2_c1 = nS_st3_b2_c1;
  assign nS_st4_b3_c1 = nS_st3_b3_c1;
  assign nS_st4_b4_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b4_c0 : nS_st3_b4_c1;
  assign nS_st4_b5_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b5_c0 : nS_st3_b5_c1;
  assign nS_st4_b6_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b6_c0 : nS_st3_b6_c1;
  assign nS_st4_b7_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b7_c0 : nS_st3_b7_c1;
  assign nS_st4_b8_c1 = nS_st3_b8_c1;
  assign nS_st4_b9_c1 = nS_st3_b9_c1;
  assign nS_st4_b10_c1 = nS_st3_b10_c1;
  assign nS_st4_b11_c1 = nS_st3_b11_c1;
  assign nS_st4_b12_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b12_c0 : nS_st3_b12_c1;
  assign nS_st4_b13_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b13_c0 : nS_st3_b13_c1;
  assign nS_st4_b14_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b14_c0 : nS_st3_b14_c1;
  assign nS_st4_b15_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b15_c0 : nS_st3_b15_c1;
  assign nS_st4_b16_c1 = nS_st3_b16_c1;
  assign nS_st4_b17_c1 = nS_st3_b17_c1;
  assign nS_st4_b18_c1 = nS_st3_b18_c1;
  assign nS_st4_b19_c1 = nS_st3_b19_c1;
  assign nS_st4_b20_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b20_c0 : nS_st3_b20_c1;
  assign nS_st4_b21_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b21_c0 : nS_st3_b21_c1;
  assign nS_st4_b22_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b22_c0 : nS_st3_b22_c1;
  assign nS_st4_b23_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b23_c0 : nS_st3_b23_c1;
  assign nS_st4_b24_c1 = nS_st3_b24_c1;
  assign nS_st4_b25_c1 = nS_st3_b25_c1;
  assign nS_st4_b26_c1 = nS_st3_b26_c1;
  assign nS_st4_b27_c1 = nS_st3_b27_c1;
  assign nS_st4_b28_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b28_c0 : nS_st3_b28_c1;
  assign nS_st4_b29_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b29_c0 : nS_st3_b29_c1;
  assign nS_st4_b30_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b30_c0 : nS_st3_b30_c1;
  assign nS_st4_b31_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b31_c0 : nS_st3_b31_c1;
  assign nS_st4_b32_c1 = nS_st3_b32_c1;
  assign nS_st4_b33_c1 = nS_st3_b33_c1;
  assign nS_st4_b34_c1 = nS_st3_b34_c1;
  assign nS_st4_b35_c1 = nS_st3_b35_c1;
  assign nS_st4_b36_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b36_c0 : nS_st3_b36_c1;
  assign nS_st4_b37_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b37_c0 : nS_st3_b37_c1;
  assign nS_st4_b38_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b38_c0 : nS_st3_b38_c1;
  assign nS_st4_b39_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b39_c0 : nS_st3_b39_c1;
  assign nS_st4_b40_c1 = nS_st3_b40_c1;
  assign nS_st4_b41_c1 = nS_st3_b41_c1;
  assign nS_st4_b42_c1 = nS_st3_b42_c1;
  assign nS_st4_b43_c1 = nS_st3_b43_c1;
  assign nS_st4_b44_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b44_c0 : nS_st3_b44_c1;
  assign nS_st4_b45_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b45_c0 : nS_st3_b45_c1;
  assign nS_st4_b46_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b46_c0 : nS_st3_b46_c1;
  assign nS_st4_b47_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b47_c0 : nS_st3_b47_c1;
  assign nS_st4_b48_c1 = nS_st3_b48_c1;
  assign nS_st4_b49_c1 = nS_st3_b49_c1;
  assign nS_st4_b50_c1 = nS_st3_b50_c1;
  assign nS_st4_b51_c1 = nS_st3_b51_c1;
  assign nS_st4_b52_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b52_c0 : nS_st3_b52_c1;
  assign nS_st4_b53_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b53_c0 : nS_st3_b53_c1;
  assign nS_st4_b54_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b54_c0 : nS_st3_b54_c1;
  assign nS_st4_b55_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b55_c0 : nS_st3_b55_c1;
  assign nS_st4_b56_c1 = nS_st3_b56_c1;
  assign nS_st4_b57_c1 = nS_st3_b57_c1;
  assign nS_st4_b58_c1 = nS_st3_b58_c1;
  assign nS_st4_b59_c1 = nS_st3_b59_c1;
  assign nS_st4_b60_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b60_c0 : nS_st3_b60_c1;
  assign nS_st4_b61_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b61_c0 : nS_st3_b61_c1;
  assign nS_st4_b62_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b62_c0 : nS_st3_b62_c1;
  assign nS_st4_b63_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b63_c0 : nS_st3_b63_c1;
  assign nS_st4_b64_c1 = nS_st3_b64_c1;
  assign nS_st4_b65_c1 = nS_st3_b65_c1;
  assign nS_st4_b66_c1 = nS_st3_b66_c1;
  assign nS_st4_b67_c1 = nS_st3_b67_c1;
  assign nS_st4_b68_c1 = (nC_st3_b67_c1 == 0) ? nS_st3_b68_c0 : nS_st3_b68_c1;
  assign nS_st4_b69_c1 = (nC_st3_b67_c1 == 0) ? nS_st3_b69_c0 : nS_st3_b69_c1;
  assign nS_st4_b70_c1 = (nC_st3_b67_c1 == 0) ? nS_st3_b70_c0 : nS_st3_b70_c1;
  assign nS_st4_b71_c1 = (nC_st3_b67_c1 == 0) ? nS_st3_b71_c0 : nS_st3_b71_c1;
  assign nS_st4_b72_c1 = nS_st3_b72_c1;
  assign nS_st4_b73_c1 = nS_st3_b73_c1;
  assign nS_st4_b74_c1 = nS_st3_b74_c1;
  assign nS_st4_b75_c1 = nS_st3_b75_c1;
  assign nS_st4_b76_c1 = (nC_st3_b75_c1 == 0) ? nS_st3_b76_c0 : nS_st3_b76_c1;
  assign nS_st4_b77_c1 = (nC_st3_b75_c1 == 0) ? nS_st3_b77_c0 : nS_st3_b77_c1;
  assign nS_st4_b78_c1 = (nC_st3_b75_c1 == 0) ? nS_st3_b78_c0 : nS_st3_b78_c1;
  assign nS_st4_b79_c1 = (nC_st3_b75_c1 == 0) ? nS_st3_b79_c0 : nS_st3_b79_c1;
  assign nS_st4_b80_c1 = nS_st3_b80_c1;
  assign nS_st4_b81_c1 = nS_st3_b81_c1;
  assign nS_st4_b82_c1 = nS_st3_b82_c1;
  assign nS_st4_b83_c1 = nS_st3_b83_c1;
  assign nS_st4_b84_c1 = (nC_st3_b83_c1 == 0) ? nS_st3_b84_c0 : nS_st3_b84_c1;
  assign nS_st4_b85_c1 = (nC_st3_b83_c1 == 0) ? nS_st3_b85_c0 : nS_st3_b85_c1;
  assign nS_st4_b86_c1 = (nC_st3_b83_c1 == 0) ? nS_st3_b86_c0 : nS_st3_b86_c1;
  assign nS_st4_b87_c1 = (nC_st3_b83_c1 == 0) ? nS_st3_b87_c0 : nS_st3_b87_c1;
  assign nS_st4_b88_c1 = nS_st3_b88_c1;
  assign nS_st4_b89_c1 = nS_st3_b89_c1;
  assign nS_st4_b90_c1 = nS_st3_b90_c1;
  assign nS_st4_b91_c1 = nS_st3_b91_c1;
  assign nS_st4_b92_c1 = (nC_st3_b91_c1 == 0) ? nS_st3_b92_c0 : nS_st3_b92_c1;
  assign nS_st4_b93_c1 = (nC_st3_b91_c1 == 0) ? nS_st3_b93_c0 : nS_st3_b93_c1;
  assign nS_st4_b94_c1 = (nC_st3_b91_c1 == 0) ? nS_st3_b94_c0 : nS_st3_b94_c1;
  assign nS_st4_b95_c1 = (nC_st3_b91_c1 == 0) ? nS_st3_b95_c0 : nS_st3_b95_c1;
  assign nS_st4_b96_c1 = nS_st3_b96_c1;
  assign nS_st4_b97_c1 = nS_st3_b97_c1;
  assign nS_st4_b98_c1 = nS_st3_b98_c1;
  assign nS_st4_b99_c1 = nS_st3_b99_c1;
  assign nS_st4_b100_c1 = (nC_st3_b99_c1 == 0) ? nS_st3_b100_c0 : nS_st3_b100_c1;
  assign nS_st4_b101_c1 = (nC_st3_b99_c1 == 0) ? nS_st3_b101_c0 : nS_st3_b101_c1;
  assign nS_st4_b102_c1 = (nC_st3_b99_c1 == 0) ? nS_st3_b102_c0 : nS_st3_b102_c1;
  assign nS_st4_b103_c1 = (nC_st3_b99_c1 == 0) ? nS_st3_b103_c0 : nS_st3_b103_c1;
  assign nS_st4_b104_c1 = nS_st3_b104_c1;
  assign nS_st4_b105_c1 = nS_st3_b105_c1;
  assign nS_st4_b106_c1 = nS_st3_b106_c1;
  assign nS_st4_b107_c1 = nS_st3_b107_c1;
  assign nS_st4_b108_c1 = (nC_st3_b107_c1 == 0) ? nS_st3_b108_c0 : nS_st3_b108_c1;
  assign nS_st4_b109_c1 = (nC_st3_b107_c1 == 0) ? nS_st3_b109_c0 : nS_st3_b109_c1;
  assign nS_st4_b110_c1 = (nC_st3_b107_c1 == 0) ? nS_st3_b110_c0 : nS_st3_b110_c1;
  assign nS_st4_b111_c1 = (nC_st3_b107_c1 == 0) ? nS_st3_b111_c0 : nS_st3_b111_c1;
  assign nS_st4_b112_c1 = nS_st3_b112_c1;
  assign nS_st4_b113_c1 = nS_st3_b113_c1;
  assign nS_st4_b114_c1 = nS_st3_b114_c1;
  assign nS_st4_b115_c1 = nS_st3_b115_c1;
  assign nS_st4_b116_c1 = (nC_st3_b115_c1 == 0) ? nS_st3_b116_c0 : nS_st3_b116_c1;
  assign nS_st4_b117_c1 = (nC_st3_b115_c1 == 0) ? nS_st3_b117_c0 : nS_st3_b117_c1;
  assign nS_st4_b118_c1 = (nC_st3_b115_c1 == 0) ? nS_st3_b118_c0 : nS_st3_b118_c1;
  assign nS_st4_b119_c1 = (nC_st3_b115_c1 == 0) ? nS_st3_b119_c0 : nS_st3_b119_c1;
  assign nS_st4_b120_c1 = nS_st3_b120_c1;
  assign nS_st4_b121_c1 = nS_st3_b121_c1;
  assign nS_st4_b122_c1 = nS_st3_b122_c1;
  assign nS_st4_b123_c1 = nS_st3_b123_c1;
  assign nS_st4_b124_c1 = (nC_st3_b123_c1 == 0) ? nS_st3_b124_c0 : nS_st3_b124_c1;
  assign nS_st4_b125_c1 = (nC_st3_b123_c1 == 0) ? nS_st3_b125_c0 : nS_st3_b125_c1;
  assign nS_st4_b126_c1 = (nC_st3_b123_c1 == 0) ? nS_st3_b126_c0 : nS_st3_b126_c1;
  assign nS_st4_b127_c1 = (nC_st3_b123_c1 == 0) ? nS_st3_b127_c0 : nS_st3_b127_c1;
  assign nS_st4_b128_c1 = nS_st3_b128_c1;
  assign nS_st4_b129_c1 = nS_st3_b129_c1;
  assign nS_st4_b130_c1 = nS_st3_b130_c1;
  assign nS_st4_b131_c1 = nS_st3_b131_c1;
  assign nS_st4_b132_c1 = (nC_st3_b131_c1 == 0) ? nS_st3_b132_c0 : nS_st3_b132_c1;
  assign nS_st4_b133_c1 = (nC_st3_b131_c1 == 0) ? nS_st3_b133_c0 : nS_st3_b133_c1;
  assign nS_st4_b134_c1 = (nC_st3_b131_c1 == 0) ? nS_st3_b134_c0 : nS_st3_b134_c1;
  assign nS_st4_b135_c1 = (nC_st3_b131_c1 == 0) ? nS_st3_b135_c0 : nS_st3_b135_c1;
  assign nS_st4_b136_c1 = nS_st3_b136_c1;
  assign nS_st4_b137_c1 = nS_st3_b137_c1;
  assign nS_st4_b138_c1 = nS_st3_b138_c1;
  assign nS_st4_b139_c1 = nS_st3_b139_c1;
  assign nS_st4_b140_c1 = (nC_st3_b139_c1 == 0) ? nS_st3_b140_c0 : nS_st3_b140_c1;
  assign nS_st4_b141_c1 = (nC_st3_b139_c1 == 0) ? nS_st3_b141_c0 : nS_st3_b141_c1;
  assign nS_st4_b142_c1 = (nC_st3_b139_c1 == 0) ? nS_st3_b142_c0 : nS_st3_b142_c1;
  assign nS_st4_b143_c1 = (nC_st3_b139_c1 == 0) ? nS_st3_b143_c0 : nS_st3_b143_c1;
  assign nS_st4_b144_c1 = nS_st3_b144_c1;
  assign nS_st4_b145_c1 = nS_st3_b145_c1;
  assign nS_st4_b146_c1 = nS_st3_b146_c1;
  assign nS_st4_b147_c1 = nS_st3_b147_c1;
  assign nS_st4_b148_c1 = (nC_st3_b147_c1 == 0) ? nS_st3_b148_c0 : nS_st3_b148_c1;
  assign nS_st4_b149_c1 = (nC_st3_b147_c1 == 0) ? nS_st3_b149_c0 : nS_st3_b149_c1;
  assign nS_st4_b150_c1 = (nC_st3_b147_c1 == 0) ? nS_st3_b150_c0 : nS_st3_b150_c1;
  assign nS_st4_b151_c1 = (nC_st3_b147_c1 == 0) ? nS_st3_b151_c0 : nS_st3_b151_c1;
  assign nS_st4_b152_c1 = nS_st3_b152_c1;
  assign nS_st4_b153_c1 = nS_st3_b153_c1;
  assign nS_st4_b154_c1 = nS_st3_b154_c1;
  assign nS_st4_b155_c1 = nS_st3_b155_c1;
  assign nS_st4_b156_c1 = (nC_st3_b155_c1 == 0) ? nS_st3_b156_c0 : nS_st3_b156_c1;
  assign nS_st4_b157_c1 = (nC_st3_b155_c1 == 0) ? nS_st3_b157_c0 : nS_st3_b157_c1;
  assign nS_st4_b158_c1 = (nC_st3_b155_c1 == 0) ? nS_st3_b158_c0 : nS_st3_b158_c1;
  assign nS_st4_b159_c1 = (nC_st3_b155_c1 == 0) ? nS_st3_b159_c0 : nS_st3_b159_c1;
  assign nS_st4_b160_c1 = nS_st3_b160_c1;
  assign nS_st4_b161_c1 = nS_st3_b161_c1;
  assign nS_st4_b162_c1 = nS_st3_b162_c1;
  assign nS_st4_b163_c1 = nS_st3_b163_c1;
  assign nS_st4_b164_c1 = (nC_st3_b163_c1 == 0) ? nS_st3_b164_c0 : nS_st3_b164_c1;
  assign nS_st4_b165_c1 = (nC_st3_b163_c1 == 0) ? nS_st3_b165_c0 : nS_st3_b165_c1;
  assign nS_st4_b166_c1 = (nC_st3_b163_c1 == 0) ? nS_st3_b166_c0 : nS_st3_b166_c1;
  assign nS_st4_b167_c1 = (nC_st3_b163_c1 == 0) ? nS_st3_b167_c0 : nS_st3_b167_c1;
  assign nS_st4_b168_c1 = nS_st3_b168_c1;
  assign nS_st4_b169_c1 = nS_st3_b169_c1;
  assign nS_st4_b170_c1 = nS_st3_b170_c1;
  assign nS_st4_b171_c1 = nS_st3_b171_c1;
  assign nS_st4_b172_c1 = (nC_st3_b171_c1 == 0) ? nS_st3_b172_c0 : nS_st3_b172_c1;
  assign nS_st4_b173_c1 = (nC_st3_b171_c1 == 0) ? nS_st3_b173_c0 : nS_st3_b173_c1;
  assign nS_st4_b174_c1 = (nC_st3_b171_c1 == 0) ? nS_st3_b174_c0 : nS_st3_b174_c1;
  assign nS_st4_b175_c1 = (nC_st3_b171_c1 == 0) ? nS_st3_b175_c0 : nS_st3_b175_c1;
  assign nS_st4_b176_c1 = nS_st3_b176_c1;
  assign nS_st4_b177_c1 = nS_st3_b177_c1;
  assign nS_st4_b178_c1 = nS_st3_b178_c1;
  assign nS_st4_b179_c1 = nS_st3_b179_c1;
  assign nS_st4_b180_c1 = (nC_st3_b179_c1 == 0) ? nS_st3_b180_c0 : nS_st3_b180_c1;
  assign nS_st4_b181_c1 = (nC_st3_b179_c1 == 0) ? nS_st3_b181_c0 : nS_st3_b181_c1;
  assign nS_st4_b182_c1 = (nC_st3_b179_c1 == 0) ? nS_st3_b182_c0 : nS_st3_b182_c1;
  assign nS_st4_b183_c1 = (nC_st3_b179_c1 == 0) ? nS_st3_b183_c0 : nS_st3_b183_c1;
  assign nS_st4_b184_c1 = nS_st3_b184_c1;
  assign nS_st4_b185_c1 = nS_st3_b185_c1;
  assign nS_st4_b186_c1 = nS_st3_b186_c1;
  assign nS_st4_b187_c1 = nS_st3_b187_c1;
  assign nS_st4_b188_c1 = (nC_st3_b187_c1 == 0) ? nS_st3_b188_c0 : nS_st3_b188_c1;
  assign nS_st4_b189_c1 = (nC_st3_b187_c1 == 0) ? nS_st3_b189_c0 : nS_st3_b189_c1;
  assign nS_st4_b190_c1 = (nC_st3_b187_c1 == 0) ? nS_st3_b190_c0 : nS_st3_b190_c1;
  assign nS_st4_b191_c1 = (nC_st3_b187_c1 == 0) ? nS_st3_b191_c0 : nS_st3_b191_c1;
  assign nS_st4_b192_c1 = nS_st3_b192_c1;
  assign nS_st4_b193_c1 = nS_st3_b193_c1;
  assign nS_st4_b194_c1 = nS_st3_b194_c1;
  assign nS_st4_b195_c1 = nS_st3_b195_c1;
  assign nS_st4_b196_c1 = (nC_st3_b195_c1 == 0) ? nS_st3_b196_c0 : nS_st3_b196_c1;
  assign nS_st4_b197_c1 = (nC_st3_b195_c1 == 0) ? nS_st3_b197_c0 : nS_st3_b197_c1;
  assign nS_st4_b198_c1 = (nC_st3_b195_c1 == 0) ? nS_st3_b198_c0 : nS_st3_b198_c1;
  assign nS_st4_b199_c1 = (nC_st3_b195_c1 == 0) ? nS_st3_b199_c0 : nS_st3_b199_c1;
  assign nS_st4_b200_c1 = nS_st3_b200_c1;
  assign nS_st4_b201_c1 = nS_st3_b201_c1;
  assign nS_st4_b202_c1 = nS_st3_b202_c1;
  assign nS_st4_b203_c1 = nS_st3_b203_c1;
  assign nS_st4_b204_c1 = (nC_st3_b203_c1 == 0) ? nS_st3_b204_c0 : nS_st3_b204_c1;
  assign nS_st4_b205_c1 = (nC_st3_b203_c1 == 0) ? nS_st3_b205_c0 : nS_st3_b205_c1;
  assign nS_st4_b206_c1 = (nC_st3_b203_c1 == 0) ? nS_st3_b206_c0 : nS_st3_b206_c1;
  assign nS_st4_b207_c1 = (nC_st3_b203_c1 == 0) ? nS_st3_b207_c0 : nS_st3_b207_c1;
  assign nS_st4_b208_c1 = nS_st3_b208_c1;
  assign nS_st4_b209_c1 = nS_st3_b209_c1;
  assign nS_st4_b210_c1 = nS_st3_b210_c1;
  assign nS_st4_b211_c1 = nS_st3_b211_c1;
  assign nS_st4_b212_c1 = (nC_st3_b211_c1 == 0) ? nS_st3_b212_c0 : nS_st3_b212_c1;
  assign nS_st4_b213_c1 = (nC_st3_b211_c1 == 0) ? nS_st3_b213_c0 : nS_st3_b213_c1;
  assign nS_st4_b214_c1 = (nC_st3_b211_c1 == 0) ? nS_st3_b214_c0 : nS_st3_b214_c1;
  assign nS_st4_b215_c1 = (nC_st3_b211_c1 == 0) ? nS_st3_b215_c0 : nS_st3_b215_c1;
  assign nS_st4_b216_c1 = nS_st3_b216_c1;
  assign nS_st4_b217_c1 = nS_st3_b217_c1;
  assign nS_st4_b218_c1 = nS_st3_b218_c1;
  assign nS_st4_b219_c1 = nS_st3_b219_c1;
  assign nS_st4_b220_c1 = (nC_st3_b219_c1 == 0) ? nS_st3_b220_c0 : nS_st3_b220_c1;
  assign nS_st4_b221_c1 = (nC_st3_b219_c1 == 0) ? nS_st3_b221_c0 : nS_st3_b221_c1;
  assign nS_st4_b222_c1 = (nC_st3_b219_c1 == 0) ? nS_st3_b222_c0 : nS_st3_b222_c1;
  assign nS_st4_b223_c1 = (nC_st3_b219_c1 == 0) ? nS_st3_b223_c0 : nS_st3_b223_c1;
  assign nS_st4_b224_c1 = nS_st3_b224_c1;
  assign nS_st4_b225_c1 = nS_st3_b225_c1;
  assign nS_st4_b226_c1 = nS_st3_b226_c1;
  assign nS_st4_b227_c1 = nS_st3_b227_c1;
  assign nS_st4_b228_c1 = (nC_st3_b227_c1 == 0) ? nS_st3_b228_c0 : nS_st3_b228_c1;
  assign nS_st4_b229_c1 = (nC_st3_b227_c1 == 0) ? nS_st3_b229_c0 : nS_st3_b229_c1;
  assign nS_st4_b230_c1 = (nC_st3_b227_c1 == 0) ? nS_st3_b230_c0 : nS_st3_b230_c1;
  assign nS_st4_b231_c1 = (nC_st3_b227_c1 == 0) ? nS_st3_b231_c0 : nS_st3_b231_c1;
  assign nS_st4_b232_c1 = nS_st3_b232_c1;
  assign nS_st4_b233_c1 = nS_st3_b233_c1;
  assign nS_st4_b234_c1 = nS_st3_b234_c1;
  assign nS_st4_b235_c1 = nS_st3_b235_c1;
  assign nS_st4_b236_c1 = (nC_st3_b235_c1 == 0) ? nS_st3_b236_c0 : nS_st3_b236_c1;
  assign nS_st4_b237_c1 = (nC_st3_b235_c1 == 0) ? nS_st3_b237_c0 : nS_st3_b237_c1;
  assign nS_st4_b238_c1 = (nC_st3_b235_c1 == 0) ? nS_st3_b238_c0 : nS_st3_b238_c1;
  assign nS_st4_b239_c1 = (nC_st3_b235_c1 == 0) ? nS_st3_b239_c0 : nS_st3_b239_c1;
  assign nS_st4_b240_c1 = nS_st3_b240_c1;
  assign nS_st4_b241_c1 = nS_st3_b241_c1;
  assign nS_st4_b242_c1 = nS_st3_b242_c1;
  assign nS_st4_b243_c1 = nS_st3_b243_c1;
  assign nS_st4_b244_c1 = (nC_st3_b243_c1 == 0) ? nS_st3_b244_c0 : nS_st3_b244_c1;
  assign nS_st4_b245_c1 = (nC_st3_b243_c1 == 0) ? nS_st3_b245_c0 : nS_st3_b245_c1;
  assign nS_st4_b246_c1 = (nC_st3_b243_c1 == 0) ? nS_st3_b246_c0 : nS_st3_b246_c1;
  assign nS_st4_b247_c1 = (nC_st3_b243_c1 == 0) ? nS_st3_b247_c0 : nS_st3_b247_c1;
  assign nS_st4_b248_c1 = nS_st3_b248_c1;
  assign nS_st4_b249_c1 = nS_st3_b249_c1;
  assign nS_st4_b250_c1 = nS_st3_b250_c1;
  assign nS_st4_b251_c1 = nS_st3_b251_c1;
  assign nS_st4_b252_c1 = (nC_st3_b251_c1 == 0) ? nS_st3_b252_c0 : nS_st3_b252_c1;
  assign nS_st4_b253_c1 = (nC_st3_b251_c1 == 0) ? nS_st3_b253_c0 : nS_st3_b253_c1;
  assign nS_st4_b254_c1 = (nC_st3_b251_c1 == 0) ? nS_st3_b254_c0 : nS_st3_b254_c1;
  assign nS_st4_b255_c1 = (nC_st3_b251_c1 == 0) ? nS_st3_b255_c0 : nS_st3_b255_c1;
  assign nC_st4_b7_c0 = (nC_st3_b3_c0 == 0) ? nC_st3_b7_c0 : nC_st3_b7_c1;
  assign nC_st4_b15_c0 = (nC_st3_b11_c0 == 0) ? nC_st3_b15_c0 : nC_st3_b15_c1;
  assign nC_st4_b23_c0 = (nC_st3_b19_c0 == 0) ? nC_st3_b23_c0 : nC_st3_b23_c1;
  assign nC_st4_b31_c0 = (nC_st3_b27_c0 == 0) ? nC_st3_b31_c0 : nC_st3_b31_c1;
  assign nC_st4_b39_c0 = (nC_st3_b35_c0 == 0) ? nC_st3_b39_c0 : nC_st3_b39_c1;
  assign nC_st4_b47_c0 = (nC_st3_b43_c0 == 0) ? nC_st3_b47_c0 : nC_st3_b47_c1;
  assign nC_st4_b55_c0 = (nC_st3_b51_c0 == 0) ? nC_st3_b55_c0 : nC_st3_b55_c1;
  assign nC_st4_b63_c0 = (nC_st3_b59_c0 == 0) ? nC_st3_b63_c0 : nC_st3_b63_c1;
  assign nC_st4_b71_c0 = (nC_st3_b67_c0 == 0) ? nC_st3_b71_c0 : nC_st3_b71_c1;
  assign nC_st4_b79_c0 = (nC_st3_b75_c0 == 0) ? nC_st3_b79_c0 : nC_st3_b79_c1;
  assign nC_st4_b87_c0 = (nC_st3_b83_c0 == 0) ? nC_st3_b87_c0 : nC_st3_b87_c1;
  assign nC_st4_b95_c0 = (nC_st3_b91_c0 == 0) ? nC_st3_b95_c0 : nC_st3_b95_c1;
  assign nC_st4_b103_c0 = (nC_st3_b99_c0 == 0) ? nC_st3_b103_c0 : nC_st3_b103_c1;
  assign nC_st4_b111_c0 = (nC_st3_b107_c0 == 0) ? nC_st3_b111_c0 : nC_st3_b111_c1;
  assign nC_st4_b119_c0 = (nC_st3_b115_c0 == 0) ? nC_st3_b119_c0 : nC_st3_b119_c1;
  assign nC_st4_b127_c0 = (nC_st3_b123_c0 == 0) ? nC_st3_b127_c0 : nC_st3_b127_c1;
  assign nC_st4_b135_c0 = (nC_st3_b131_c0 == 0) ? nC_st3_b135_c0 : nC_st3_b135_c1;
  assign nC_st4_b143_c0 = (nC_st3_b139_c0 == 0) ? nC_st3_b143_c0 : nC_st3_b143_c1;
  assign nC_st4_b151_c0 = (nC_st3_b147_c0 == 0) ? nC_st3_b151_c0 : nC_st3_b151_c1;
  assign nC_st4_b159_c0 = (nC_st3_b155_c0 == 0) ? nC_st3_b159_c0 : nC_st3_b159_c1;
  assign nC_st4_b167_c0 = (nC_st3_b163_c0 == 0) ? nC_st3_b167_c0 : nC_st3_b167_c1;
  assign nC_st4_b175_c0 = (nC_st3_b171_c0 == 0) ? nC_st3_b175_c0 : nC_st3_b175_c1;
  assign nC_st4_b183_c0 = (nC_st3_b179_c0 == 0) ? nC_st3_b183_c0 : nC_st3_b183_c1;
  assign nC_st4_b191_c0 = (nC_st3_b187_c0 == 0) ? nC_st3_b191_c0 : nC_st3_b191_c1;
  assign nC_st4_b199_c0 = (nC_st3_b195_c0 == 0) ? nC_st3_b199_c0 : nC_st3_b199_c1;
  assign nC_st4_b207_c0 = (nC_st3_b203_c0 == 0) ? nC_st3_b207_c0 : nC_st3_b207_c1;
  assign nC_st4_b215_c0 = (nC_st3_b211_c0 == 0) ? nC_st3_b215_c0 : nC_st3_b215_c1;
  assign nC_st4_b223_c0 = (nC_st3_b219_c0 == 0) ? nC_st3_b223_c0 : nC_st3_b223_c1;
  assign nC_st4_b231_c0 = (nC_st3_b227_c0 == 0) ? nC_st3_b231_c0 : nC_st3_b231_c1;
  assign nC_st4_b239_c0 = (nC_st3_b235_c0 == 0) ? nC_st3_b239_c0 : nC_st3_b239_c1;
  assign nC_st4_b247_c0 = (nC_st3_b243_c0 == 0) ? nC_st3_b247_c0 : nC_st3_b247_c1;
  assign nC_st4_b255_c0 = (nC_st3_b251_c0 == 0) ? nC_st3_b255_c0 : nC_st3_b255_c1;
  assign nC_st4_b7_c1 = (nC_st3_b3_c1 == 0) ? nC_st3_b7_c0 : nC_st3_b7_c1;
  assign nC_st4_b15_c1 = (nC_st3_b11_c1 == 0) ? nC_st3_b15_c0 : nC_st3_b15_c1;
  assign nC_st4_b23_c1 = (nC_st3_b19_c1 == 0) ? nC_st3_b23_c0 : nC_st3_b23_c1;
  assign nC_st4_b31_c1 = (nC_st3_b27_c1 == 0) ? nC_st3_b31_c0 : nC_st3_b31_c1;
  assign nC_st4_b39_c1 = (nC_st3_b35_c1 == 0) ? nC_st3_b39_c0 : nC_st3_b39_c1;
  assign nC_st4_b47_c1 = (nC_st3_b43_c1 == 0) ? nC_st3_b47_c0 : nC_st3_b47_c1;
  assign nC_st4_b55_c1 = (nC_st3_b51_c1 == 0) ? nC_st3_b55_c0 : nC_st3_b55_c1;
  assign nC_st4_b63_c1 = (nC_st3_b59_c1 == 0) ? nC_st3_b63_c0 : nC_st3_b63_c1;
  assign nC_st4_b71_c1 = (nC_st3_b67_c1 == 0) ? nC_st3_b71_c0 : nC_st3_b71_c1;
  assign nC_st4_b79_c1 = (nC_st3_b75_c1 == 0) ? nC_st3_b79_c0 : nC_st3_b79_c1;
  assign nC_st4_b87_c1 = (nC_st3_b83_c1 == 0) ? nC_st3_b87_c0 : nC_st3_b87_c1;
  assign nC_st4_b95_c1 = (nC_st3_b91_c1 == 0) ? nC_st3_b95_c0 : nC_st3_b95_c1;
  assign nC_st4_b103_c1 = (nC_st3_b99_c1 == 0) ? nC_st3_b103_c0 : nC_st3_b103_c1;
  assign nC_st4_b111_c1 = (nC_st3_b107_c1 == 0) ? nC_st3_b111_c0 : nC_st3_b111_c1;
  assign nC_st4_b119_c1 = (nC_st3_b115_c1 == 0) ? nC_st3_b119_c0 : nC_st3_b119_c1;
  assign nC_st4_b127_c1 = (nC_st3_b123_c1 == 0) ? nC_st3_b127_c0 : nC_st3_b127_c1;
  assign nC_st4_b135_c1 = (nC_st3_b131_c1 == 0) ? nC_st3_b135_c0 : nC_st3_b135_c1;
  assign nC_st4_b143_c1 = (nC_st3_b139_c1 == 0) ? nC_st3_b143_c0 : nC_st3_b143_c1;
  assign nC_st4_b151_c1 = (nC_st3_b147_c1 == 0) ? nC_st3_b151_c0 : nC_st3_b151_c1;
  assign nC_st4_b159_c1 = (nC_st3_b155_c1 == 0) ? nC_st3_b159_c0 : nC_st3_b159_c1;
  assign nC_st4_b167_c1 = (nC_st3_b163_c1 == 0) ? nC_st3_b167_c0 : nC_st3_b167_c1;
  assign nC_st4_b175_c1 = (nC_st3_b171_c1 == 0) ? nC_st3_b175_c0 : nC_st3_b175_c1;
  assign nC_st4_b183_c1 = (nC_st3_b179_c1 == 0) ? nC_st3_b183_c0 : nC_st3_b183_c1;
  assign nC_st4_b191_c1 = (nC_st3_b187_c1 == 0) ? nC_st3_b191_c0 : nC_st3_b191_c1;
  assign nC_st4_b199_c1 = (nC_st3_b195_c1 == 0) ? nC_st3_b199_c0 : nC_st3_b199_c1;
  assign nC_st4_b207_c1 = (nC_st3_b203_c1 == 0) ? nC_st3_b207_c0 : nC_st3_b207_c1;
  assign nC_st4_b215_c1 = (nC_st3_b211_c1 == 0) ? nC_st3_b215_c0 : nC_st3_b215_c1;
  assign nC_st4_b223_c1 = (nC_st3_b219_c1 == 0) ? nC_st3_b223_c0 : nC_st3_b223_c1;
  assign nC_st4_b231_c1 = (nC_st3_b227_c1 == 0) ? nC_st3_b231_c0 : nC_st3_b231_c1;
  assign nC_st4_b239_c1 = (nC_st3_b235_c1 == 0) ? nC_st3_b239_c0 : nC_st3_b239_c1;
  assign nC_st4_b247_c1 = (nC_st3_b243_c1 == 0) ? nC_st3_b247_c0 : nC_st3_b247_c1;
  assign nC_st4_b255_c1 = (nC_st3_b251_c1 == 0) ? nC_st3_b255_c0 : nC_st3_b255_c1;

  assign nS_st5_b0_c0 = nS_st4_b0_c0;
  assign nS_st5_b1_c0 = nS_st4_b1_c0;
  assign nS_st5_b2_c0 = nS_st4_b2_c0;
  assign nS_st5_b3_c0 = nS_st4_b3_c0;
  assign nS_st5_b4_c0 = nS_st4_b4_c0;
  assign nS_st5_b5_c0 = nS_st4_b5_c0;
  assign nS_st5_b6_c0 = nS_st4_b6_c0;
  assign nS_st5_b7_c0 = nS_st4_b7_c0;
  assign nS_st5_b8_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b8_c0 : nS_st4_b8_c1;
  assign nS_st5_b9_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b9_c0 : nS_st4_b9_c1;
  assign nS_st5_b10_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b10_c0 : nS_st4_b10_c1;
  assign nS_st5_b11_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b11_c0 : nS_st4_b11_c1;
  assign nS_st5_b12_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b12_c0 : nS_st4_b12_c1;
  assign nS_st5_b13_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b13_c0 : nS_st4_b13_c1;
  assign nS_st5_b14_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b14_c0 : nS_st4_b14_c1;
  assign nS_st5_b15_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b15_c0 : nS_st4_b15_c1;
  assign nS_st5_b16_c0 = nS_st4_b16_c0;
  assign nS_st5_b17_c0 = nS_st4_b17_c0;
  assign nS_st5_b18_c0 = nS_st4_b18_c0;
  assign nS_st5_b19_c0 = nS_st4_b19_c0;
  assign nS_st5_b20_c0 = nS_st4_b20_c0;
  assign nS_st5_b21_c0 = nS_st4_b21_c0;
  assign nS_st5_b22_c0 = nS_st4_b22_c0;
  assign nS_st5_b23_c0 = nS_st4_b23_c0;
  assign nS_st5_b24_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b24_c0 : nS_st4_b24_c1;
  assign nS_st5_b25_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b25_c0 : nS_st4_b25_c1;
  assign nS_st5_b26_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b26_c0 : nS_st4_b26_c1;
  assign nS_st5_b27_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b27_c0 : nS_st4_b27_c1;
  assign nS_st5_b28_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b28_c0 : nS_st4_b28_c1;
  assign nS_st5_b29_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b29_c0 : nS_st4_b29_c1;
  assign nS_st5_b30_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b30_c0 : nS_st4_b30_c1;
  assign nS_st5_b31_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b31_c0 : nS_st4_b31_c1;
  assign nS_st5_b32_c0 = nS_st4_b32_c0;
  assign nS_st5_b33_c0 = nS_st4_b33_c0;
  assign nS_st5_b34_c0 = nS_st4_b34_c0;
  assign nS_st5_b35_c0 = nS_st4_b35_c0;
  assign nS_st5_b36_c0 = nS_st4_b36_c0;
  assign nS_st5_b37_c0 = nS_st4_b37_c0;
  assign nS_st5_b38_c0 = nS_st4_b38_c0;
  assign nS_st5_b39_c0 = nS_st4_b39_c0;
  assign nS_st5_b40_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b40_c0 : nS_st4_b40_c1;
  assign nS_st5_b41_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b41_c0 : nS_st4_b41_c1;
  assign nS_st5_b42_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b42_c0 : nS_st4_b42_c1;
  assign nS_st5_b43_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b43_c0 : nS_st4_b43_c1;
  assign nS_st5_b44_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b44_c0 : nS_st4_b44_c1;
  assign nS_st5_b45_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b45_c0 : nS_st4_b45_c1;
  assign nS_st5_b46_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b46_c0 : nS_st4_b46_c1;
  assign nS_st5_b47_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b47_c0 : nS_st4_b47_c1;
  assign nS_st5_b48_c0 = nS_st4_b48_c0;
  assign nS_st5_b49_c0 = nS_st4_b49_c0;
  assign nS_st5_b50_c0 = nS_st4_b50_c0;
  assign nS_st5_b51_c0 = nS_st4_b51_c0;
  assign nS_st5_b52_c0 = nS_st4_b52_c0;
  assign nS_st5_b53_c0 = nS_st4_b53_c0;
  assign nS_st5_b54_c0 = nS_st4_b54_c0;
  assign nS_st5_b55_c0 = nS_st4_b55_c0;
  assign nS_st5_b56_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b56_c0 : nS_st4_b56_c1;
  assign nS_st5_b57_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b57_c0 : nS_st4_b57_c1;
  assign nS_st5_b58_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b58_c0 : nS_st4_b58_c1;
  assign nS_st5_b59_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b59_c0 : nS_st4_b59_c1;
  assign nS_st5_b60_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b60_c0 : nS_st4_b60_c1;
  assign nS_st5_b61_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b61_c0 : nS_st4_b61_c1;
  assign nS_st5_b62_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b62_c0 : nS_st4_b62_c1;
  assign nS_st5_b63_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b63_c0 : nS_st4_b63_c1;
  assign nS_st5_b64_c0 = nS_st4_b64_c0;
  assign nS_st5_b65_c0 = nS_st4_b65_c0;
  assign nS_st5_b66_c0 = nS_st4_b66_c0;
  assign nS_st5_b67_c0 = nS_st4_b67_c0;
  assign nS_st5_b68_c0 = nS_st4_b68_c0;
  assign nS_st5_b69_c0 = nS_st4_b69_c0;
  assign nS_st5_b70_c0 = nS_st4_b70_c0;
  assign nS_st5_b71_c0 = nS_st4_b71_c0;
  assign nS_st5_b72_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b72_c0 : nS_st4_b72_c1;
  assign nS_st5_b73_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b73_c0 : nS_st4_b73_c1;
  assign nS_st5_b74_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b74_c0 : nS_st4_b74_c1;
  assign nS_st5_b75_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b75_c0 : nS_st4_b75_c1;
  assign nS_st5_b76_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b76_c0 : nS_st4_b76_c1;
  assign nS_st5_b77_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b77_c0 : nS_st4_b77_c1;
  assign nS_st5_b78_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b78_c0 : nS_st4_b78_c1;
  assign nS_st5_b79_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b79_c0 : nS_st4_b79_c1;
  assign nS_st5_b80_c0 = nS_st4_b80_c0;
  assign nS_st5_b81_c0 = nS_st4_b81_c0;
  assign nS_st5_b82_c0 = nS_st4_b82_c0;
  assign nS_st5_b83_c0 = nS_st4_b83_c0;
  assign nS_st5_b84_c0 = nS_st4_b84_c0;
  assign nS_st5_b85_c0 = nS_st4_b85_c0;
  assign nS_st5_b86_c0 = nS_st4_b86_c0;
  assign nS_st5_b87_c0 = nS_st4_b87_c0;
  assign nS_st5_b88_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b88_c0 : nS_st4_b88_c1;
  assign nS_st5_b89_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b89_c0 : nS_st4_b89_c1;
  assign nS_st5_b90_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b90_c0 : nS_st4_b90_c1;
  assign nS_st5_b91_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b91_c0 : nS_st4_b91_c1;
  assign nS_st5_b92_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b92_c0 : nS_st4_b92_c1;
  assign nS_st5_b93_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b93_c0 : nS_st4_b93_c1;
  assign nS_st5_b94_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b94_c0 : nS_st4_b94_c1;
  assign nS_st5_b95_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b95_c0 : nS_st4_b95_c1;
  assign nS_st5_b96_c0 = nS_st4_b96_c0;
  assign nS_st5_b97_c0 = nS_st4_b97_c0;
  assign nS_st5_b98_c0 = nS_st4_b98_c0;
  assign nS_st5_b99_c0 = nS_st4_b99_c0;
  assign nS_st5_b100_c0 = nS_st4_b100_c0;
  assign nS_st5_b101_c0 = nS_st4_b101_c0;
  assign nS_st5_b102_c0 = nS_st4_b102_c0;
  assign nS_st5_b103_c0 = nS_st4_b103_c0;
  assign nS_st5_b104_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b104_c0 : nS_st4_b104_c1;
  assign nS_st5_b105_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b105_c0 : nS_st4_b105_c1;
  assign nS_st5_b106_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b106_c0 : nS_st4_b106_c1;
  assign nS_st5_b107_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b107_c0 : nS_st4_b107_c1;
  assign nS_st5_b108_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b108_c0 : nS_st4_b108_c1;
  assign nS_st5_b109_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b109_c0 : nS_st4_b109_c1;
  assign nS_st5_b110_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b110_c0 : nS_st4_b110_c1;
  assign nS_st5_b111_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b111_c0 : nS_st4_b111_c1;
  assign nS_st5_b112_c0 = nS_st4_b112_c0;
  assign nS_st5_b113_c0 = nS_st4_b113_c0;
  assign nS_st5_b114_c0 = nS_st4_b114_c0;
  assign nS_st5_b115_c0 = nS_st4_b115_c0;
  assign nS_st5_b116_c0 = nS_st4_b116_c0;
  assign nS_st5_b117_c0 = nS_st4_b117_c0;
  assign nS_st5_b118_c0 = nS_st4_b118_c0;
  assign nS_st5_b119_c0 = nS_st4_b119_c0;
  assign nS_st5_b120_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b120_c0 : nS_st4_b120_c1;
  assign nS_st5_b121_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b121_c0 : nS_st4_b121_c1;
  assign nS_st5_b122_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b122_c0 : nS_st4_b122_c1;
  assign nS_st5_b123_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b123_c0 : nS_st4_b123_c1;
  assign nS_st5_b124_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b124_c0 : nS_st4_b124_c1;
  assign nS_st5_b125_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b125_c0 : nS_st4_b125_c1;
  assign nS_st5_b126_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b126_c0 : nS_st4_b126_c1;
  assign nS_st5_b127_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b127_c0 : nS_st4_b127_c1;
  assign nS_st5_b128_c0 = nS_st4_b128_c0;
  assign nS_st5_b129_c0 = nS_st4_b129_c0;
  assign nS_st5_b130_c0 = nS_st4_b130_c0;
  assign nS_st5_b131_c0 = nS_st4_b131_c0;
  assign nS_st5_b132_c0 = nS_st4_b132_c0;
  assign nS_st5_b133_c0 = nS_st4_b133_c0;
  assign nS_st5_b134_c0 = nS_st4_b134_c0;
  assign nS_st5_b135_c0 = nS_st4_b135_c0;
  assign nS_st5_b136_c0 = (nC_st4_b135_c0 == 0) ? nS_st4_b136_c0 : nS_st4_b136_c1;
  assign nS_st5_b137_c0 = (nC_st4_b135_c0 == 0) ? nS_st4_b137_c0 : nS_st4_b137_c1;
  assign nS_st5_b138_c0 = (nC_st4_b135_c0 == 0) ? nS_st4_b138_c0 : nS_st4_b138_c1;
  assign nS_st5_b139_c0 = (nC_st4_b135_c0 == 0) ? nS_st4_b139_c0 : nS_st4_b139_c1;
  assign nS_st5_b140_c0 = (nC_st4_b135_c0 == 0) ? nS_st4_b140_c0 : nS_st4_b140_c1;
  assign nS_st5_b141_c0 = (nC_st4_b135_c0 == 0) ? nS_st4_b141_c0 : nS_st4_b141_c1;
  assign nS_st5_b142_c0 = (nC_st4_b135_c0 == 0) ? nS_st4_b142_c0 : nS_st4_b142_c1;
  assign nS_st5_b143_c0 = (nC_st4_b135_c0 == 0) ? nS_st4_b143_c0 : nS_st4_b143_c1;
  assign nS_st5_b144_c0 = nS_st4_b144_c0;
  assign nS_st5_b145_c0 = nS_st4_b145_c0;
  assign nS_st5_b146_c0 = nS_st4_b146_c0;
  assign nS_st5_b147_c0 = nS_st4_b147_c0;
  assign nS_st5_b148_c0 = nS_st4_b148_c0;
  assign nS_st5_b149_c0 = nS_st4_b149_c0;
  assign nS_st5_b150_c0 = nS_st4_b150_c0;
  assign nS_st5_b151_c0 = nS_st4_b151_c0;
  assign nS_st5_b152_c0 = (nC_st4_b151_c0 == 0) ? nS_st4_b152_c0 : nS_st4_b152_c1;
  assign nS_st5_b153_c0 = (nC_st4_b151_c0 == 0) ? nS_st4_b153_c0 : nS_st4_b153_c1;
  assign nS_st5_b154_c0 = (nC_st4_b151_c0 == 0) ? nS_st4_b154_c0 : nS_st4_b154_c1;
  assign nS_st5_b155_c0 = (nC_st4_b151_c0 == 0) ? nS_st4_b155_c0 : nS_st4_b155_c1;
  assign nS_st5_b156_c0 = (nC_st4_b151_c0 == 0) ? nS_st4_b156_c0 : nS_st4_b156_c1;
  assign nS_st5_b157_c0 = (nC_st4_b151_c0 == 0) ? nS_st4_b157_c0 : nS_st4_b157_c1;
  assign nS_st5_b158_c0 = (nC_st4_b151_c0 == 0) ? nS_st4_b158_c0 : nS_st4_b158_c1;
  assign nS_st5_b159_c0 = (nC_st4_b151_c0 == 0) ? nS_st4_b159_c0 : nS_st4_b159_c1;
  assign nS_st5_b160_c0 = nS_st4_b160_c0;
  assign nS_st5_b161_c0 = nS_st4_b161_c0;
  assign nS_st5_b162_c0 = nS_st4_b162_c0;
  assign nS_st5_b163_c0 = nS_st4_b163_c0;
  assign nS_st5_b164_c0 = nS_st4_b164_c0;
  assign nS_st5_b165_c0 = nS_st4_b165_c0;
  assign nS_st5_b166_c0 = nS_st4_b166_c0;
  assign nS_st5_b167_c0 = nS_st4_b167_c0;
  assign nS_st5_b168_c0 = (nC_st4_b167_c0 == 0) ? nS_st4_b168_c0 : nS_st4_b168_c1;
  assign nS_st5_b169_c0 = (nC_st4_b167_c0 == 0) ? nS_st4_b169_c0 : nS_st4_b169_c1;
  assign nS_st5_b170_c0 = (nC_st4_b167_c0 == 0) ? nS_st4_b170_c0 : nS_st4_b170_c1;
  assign nS_st5_b171_c0 = (nC_st4_b167_c0 == 0) ? nS_st4_b171_c0 : nS_st4_b171_c1;
  assign nS_st5_b172_c0 = (nC_st4_b167_c0 == 0) ? nS_st4_b172_c0 : nS_st4_b172_c1;
  assign nS_st5_b173_c0 = (nC_st4_b167_c0 == 0) ? nS_st4_b173_c0 : nS_st4_b173_c1;
  assign nS_st5_b174_c0 = (nC_st4_b167_c0 == 0) ? nS_st4_b174_c0 : nS_st4_b174_c1;
  assign nS_st5_b175_c0 = (nC_st4_b167_c0 == 0) ? nS_st4_b175_c0 : nS_st4_b175_c1;
  assign nS_st5_b176_c0 = nS_st4_b176_c0;
  assign nS_st5_b177_c0 = nS_st4_b177_c0;
  assign nS_st5_b178_c0 = nS_st4_b178_c0;
  assign nS_st5_b179_c0 = nS_st4_b179_c0;
  assign nS_st5_b180_c0 = nS_st4_b180_c0;
  assign nS_st5_b181_c0 = nS_st4_b181_c0;
  assign nS_st5_b182_c0 = nS_st4_b182_c0;
  assign nS_st5_b183_c0 = nS_st4_b183_c0;
  assign nS_st5_b184_c0 = (nC_st4_b183_c0 == 0) ? nS_st4_b184_c0 : nS_st4_b184_c1;
  assign nS_st5_b185_c0 = (nC_st4_b183_c0 == 0) ? nS_st4_b185_c0 : nS_st4_b185_c1;
  assign nS_st5_b186_c0 = (nC_st4_b183_c0 == 0) ? nS_st4_b186_c0 : nS_st4_b186_c1;
  assign nS_st5_b187_c0 = (nC_st4_b183_c0 == 0) ? nS_st4_b187_c0 : nS_st4_b187_c1;
  assign nS_st5_b188_c0 = (nC_st4_b183_c0 == 0) ? nS_st4_b188_c0 : nS_st4_b188_c1;
  assign nS_st5_b189_c0 = (nC_st4_b183_c0 == 0) ? nS_st4_b189_c0 : nS_st4_b189_c1;
  assign nS_st5_b190_c0 = (nC_st4_b183_c0 == 0) ? nS_st4_b190_c0 : nS_st4_b190_c1;
  assign nS_st5_b191_c0 = (nC_st4_b183_c0 == 0) ? nS_st4_b191_c0 : nS_st4_b191_c1;
  assign nS_st5_b192_c0 = nS_st4_b192_c0;
  assign nS_st5_b193_c0 = nS_st4_b193_c0;
  assign nS_st5_b194_c0 = nS_st4_b194_c0;
  assign nS_st5_b195_c0 = nS_st4_b195_c0;
  assign nS_st5_b196_c0 = nS_st4_b196_c0;
  assign nS_st5_b197_c0 = nS_st4_b197_c0;
  assign nS_st5_b198_c0 = nS_st4_b198_c0;
  assign nS_st5_b199_c0 = nS_st4_b199_c0;
  assign nS_st5_b200_c0 = (nC_st4_b199_c0 == 0) ? nS_st4_b200_c0 : nS_st4_b200_c1;
  assign nS_st5_b201_c0 = (nC_st4_b199_c0 == 0) ? nS_st4_b201_c0 : nS_st4_b201_c1;
  assign nS_st5_b202_c0 = (nC_st4_b199_c0 == 0) ? nS_st4_b202_c0 : nS_st4_b202_c1;
  assign nS_st5_b203_c0 = (nC_st4_b199_c0 == 0) ? nS_st4_b203_c0 : nS_st4_b203_c1;
  assign nS_st5_b204_c0 = (nC_st4_b199_c0 == 0) ? nS_st4_b204_c0 : nS_st4_b204_c1;
  assign nS_st5_b205_c0 = (nC_st4_b199_c0 == 0) ? nS_st4_b205_c0 : nS_st4_b205_c1;
  assign nS_st5_b206_c0 = (nC_st4_b199_c0 == 0) ? nS_st4_b206_c0 : nS_st4_b206_c1;
  assign nS_st5_b207_c0 = (nC_st4_b199_c0 == 0) ? nS_st4_b207_c0 : nS_st4_b207_c1;
  assign nS_st5_b208_c0 = nS_st4_b208_c0;
  assign nS_st5_b209_c0 = nS_st4_b209_c0;
  assign nS_st5_b210_c0 = nS_st4_b210_c0;
  assign nS_st5_b211_c0 = nS_st4_b211_c0;
  assign nS_st5_b212_c0 = nS_st4_b212_c0;
  assign nS_st5_b213_c0 = nS_st4_b213_c0;
  assign nS_st5_b214_c0 = nS_st4_b214_c0;
  assign nS_st5_b215_c0 = nS_st4_b215_c0;
  assign nS_st5_b216_c0 = (nC_st4_b215_c0 == 0) ? nS_st4_b216_c0 : nS_st4_b216_c1;
  assign nS_st5_b217_c0 = (nC_st4_b215_c0 == 0) ? nS_st4_b217_c0 : nS_st4_b217_c1;
  assign nS_st5_b218_c0 = (nC_st4_b215_c0 == 0) ? nS_st4_b218_c0 : nS_st4_b218_c1;
  assign nS_st5_b219_c0 = (nC_st4_b215_c0 == 0) ? nS_st4_b219_c0 : nS_st4_b219_c1;
  assign nS_st5_b220_c0 = (nC_st4_b215_c0 == 0) ? nS_st4_b220_c0 : nS_st4_b220_c1;
  assign nS_st5_b221_c0 = (nC_st4_b215_c0 == 0) ? nS_st4_b221_c0 : nS_st4_b221_c1;
  assign nS_st5_b222_c0 = (nC_st4_b215_c0 == 0) ? nS_st4_b222_c0 : nS_st4_b222_c1;
  assign nS_st5_b223_c0 = (nC_st4_b215_c0 == 0) ? nS_st4_b223_c0 : nS_st4_b223_c1;
  assign nS_st5_b224_c0 = nS_st4_b224_c0;
  assign nS_st5_b225_c0 = nS_st4_b225_c0;
  assign nS_st5_b226_c0 = nS_st4_b226_c0;
  assign nS_st5_b227_c0 = nS_st4_b227_c0;
  assign nS_st5_b228_c0 = nS_st4_b228_c0;
  assign nS_st5_b229_c0 = nS_st4_b229_c0;
  assign nS_st5_b230_c0 = nS_st4_b230_c0;
  assign nS_st5_b231_c0 = nS_st4_b231_c0;
  assign nS_st5_b232_c0 = (nC_st4_b231_c0 == 0) ? nS_st4_b232_c0 : nS_st4_b232_c1;
  assign nS_st5_b233_c0 = (nC_st4_b231_c0 == 0) ? nS_st4_b233_c0 : nS_st4_b233_c1;
  assign nS_st5_b234_c0 = (nC_st4_b231_c0 == 0) ? nS_st4_b234_c0 : nS_st4_b234_c1;
  assign nS_st5_b235_c0 = (nC_st4_b231_c0 == 0) ? nS_st4_b235_c0 : nS_st4_b235_c1;
  assign nS_st5_b236_c0 = (nC_st4_b231_c0 == 0) ? nS_st4_b236_c0 : nS_st4_b236_c1;
  assign nS_st5_b237_c0 = (nC_st4_b231_c0 == 0) ? nS_st4_b237_c0 : nS_st4_b237_c1;
  assign nS_st5_b238_c0 = (nC_st4_b231_c0 == 0) ? nS_st4_b238_c0 : nS_st4_b238_c1;
  assign nS_st5_b239_c0 = (nC_st4_b231_c0 == 0) ? nS_st4_b239_c0 : nS_st4_b239_c1;
  assign nS_st5_b240_c0 = nS_st4_b240_c0;
  assign nS_st5_b241_c0 = nS_st4_b241_c0;
  assign nS_st5_b242_c0 = nS_st4_b242_c0;
  assign nS_st5_b243_c0 = nS_st4_b243_c0;
  assign nS_st5_b244_c0 = nS_st4_b244_c0;
  assign nS_st5_b245_c0 = nS_st4_b245_c0;
  assign nS_st5_b246_c0 = nS_st4_b246_c0;
  assign nS_st5_b247_c0 = nS_st4_b247_c0;
  assign nS_st5_b248_c0 = (nC_st4_b247_c0 == 0) ? nS_st4_b248_c0 : nS_st4_b248_c1;
  assign nS_st5_b249_c0 = (nC_st4_b247_c0 == 0) ? nS_st4_b249_c0 : nS_st4_b249_c1;
  assign nS_st5_b250_c0 = (nC_st4_b247_c0 == 0) ? nS_st4_b250_c0 : nS_st4_b250_c1;
  assign nS_st5_b251_c0 = (nC_st4_b247_c0 == 0) ? nS_st4_b251_c0 : nS_st4_b251_c1;
  assign nS_st5_b252_c0 = (nC_st4_b247_c0 == 0) ? nS_st4_b252_c0 : nS_st4_b252_c1;
  assign nS_st5_b253_c0 = (nC_st4_b247_c0 == 0) ? nS_st4_b253_c0 : nS_st4_b253_c1;
  assign nS_st5_b254_c0 = (nC_st4_b247_c0 == 0) ? nS_st4_b254_c0 : nS_st4_b254_c1;
  assign nS_st5_b255_c0 = (nC_st4_b247_c0 == 0) ? nS_st4_b255_c0 : nS_st4_b255_c1;
  assign nS_st5_b0_c1 = nS_st4_b0_c1;
  assign nS_st5_b1_c1 = nS_st4_b1_c1;
  assign nS_st5_b2_c1 = nS_st4_b2_c1;
  assign nS_st5_b3_c1 = nS_st4_b3_c1;
  assign nS_st5_b4_c1 = nS_st4_b4_c1;
  assign nS_st5_b5_c1 = nS_st4_b5_c1;
  assign nS_st5_b6_c1 = nS_st4_b6_c1;
  assign nS_st5_b7_c1 = nS_st4_b7_c1;
  assign nS_st5_b8_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b8_c0 : nS_st4_b8_c1;
  assign nS_st5_b9_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b9_c0 : nS_st4_b9_c1;
  assign nS_st5_b10_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b10_c0 : nS_st4_b10_c1;
  assign nS_st5_b11_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b11_c0 : nS_st4_b11_c1;
  assign nS_st5_b12_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b12_c0 : nS_st4_b12_c1;
  assign nS_st5_b13_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b13_c0 : nS_st4_b13_c1;
  assign nS_st5_b14_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b14_c0 : nS_st4_b14_c1;
  assign nS_st5_b15_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b15_c0 : nS_st4_b15_c1;
  assign nS_st5_b16_c1 = nS_st4_b16_c1;
  assign nS_st5_b17_c1 = nS_st4_b17_c1;
  assign nS_st5_b18_c1 = nS_st4_b18_c1;
  assign nS_st5_b19_c1 = nS_st4_b19_c1;
  assign nS_st5_b20_c1 = nS_st4_b20_c1;
  assign nS_st5_b21_c1 = nS_st4_b21_c1;
  assign nS_st5_b22_c1 = nS_st4_b22_c1;
  assign nS_st5_b23_c1 = nS_st4_b23_c1;
  assign nS_st5_b24_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b24_c0 : nS_st4_b24_c1;
  assign nS_st5_b25_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b25_c0 : nS_st4_b25_c1;
  assign nS_st5_b26_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b26_c0 : nS_st4_b26_c1;
  assign nS_st5_b27_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b27_c0 : nS_st4_b27_c1;
  assign nS_st5_b28_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b28_c0 : nS_st4_b28_c1;
  assign nS_st5_b29_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b29_c0 : nS_st4_b29_c1;
  assign nS_st5_b30_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b30_c0 : nS_st4_b30_c1;
  assign nS_st5_b31_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b31_c0 : nS_st4_b31_c1;
  assign nS_st5_b32_c1 = nS_st4_b32_c1;
  assign nS_st5_b33_c1 = nS_st4_b33_c1;
  assign nS_st5_b34_c1 = nS_st4_b34_c1;
  assign nS_st5_b35_c1 = nS_st4_b35_c1;
  assign nS_st5_b36_c1 = nS_st4_b36_c1;
  assign nS_st5_b37_c1 = nS_st4_b37_c1;
  assign nS_st5_b38_c1 = nS_st4_b38_c1;
  assign nS_st5_b39_c1 = nS_st4_b39_c1;
  assign nS_st5_b40_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b40_c0 : nS_st4_b40_c1;
  assign nS_st5_b41_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b41_c0 : nS_st4_b41_c1;
  assign nS_st5_b42_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b42_c0 : nS_st4_b42_c1;
  assign nS_st5_b43_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b43_c0 : nS_st4_b43_c1;
  assign nS_st5_b44_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b44_c0 : nS_st4_b44_c1;
  assign nS_st5_b45_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b45_c0 : nS_st4_b45_c1;
  assign nS_st5_b46_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b46_c0 : nS_st4_b46_c1;
  assign nS_st5_b47_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b47_c0 : nS_st4_b47_c1;
  assign nS_st5_b48_c1 = nS_st4_b48_c1;
  assign nS_st5_b49_c1 = nS_st4_b49_c1;
  assign nS_st5_b50_c1 = nS_st4_b50_c1;
  assign nS_st5_b51_c1 = nS_st4_b51_c1;
  assign nS_st5_b52_c1 = nS_st4_b52_c1;
  assign nS_st5_b53_c1 = nS_st4_b53_c1;
  assign nS_st5_b54_c1 = nS_st4_b54_c1;
  assign nS_st5_b55_c1 = nS_st4_b55_c1;
  assign nS_st5_b56_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b56_c0 : nS_st4_b56_c1;
  assign nS_st5_b57_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b57_c0 : nS_st4_b57_c1;
  assign nS_st5_b58_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b58_c0 : nS_st4_b58_c1;
  assign nS_st5_b59_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b59_c0 : nS_st4_b59_c1;
  assign nS_st5_b60_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b60_c0 : nS_st4_b60_c1;
  assign nS_st5_b61_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b61_c0 : nS_st4_b61_c1;
  assign nS_st5_b62_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b62_c0 : nS_st4_b62_c1;
  assign nS_st5_b63_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b63_c0 : nS_st4_b63_c1;
  assign nS_st5_b64_c1 = nS_st4_b64_c1;
  assign nS_st5_b65_c1 = nS_st4_b65_c1;
  assign nS_st5_b66_c1 = nS_st4_b66_c1;
  assign nS_st5_b67_c1 = nS_st4_b67_c1;
  assign nS_st5_b68_c1 = nS_st4_b68_c1;
  assign nS_st5_b69_c1 = nS_st4_b69_c1;
  assign nS_st5_b70_c1 = nS_st4_b70_c1;
  assign nS_st5_b71_c1 = nS_st4_b71_c1;
  assign nS_st5_b72_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b72_c0 : nS_st4_b72_c1;
  assign nS_st5_b73_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b73_c0 : nS_st4_b73_c1;
  assign nS_st5_b74_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b74_c0 : nS_st4_b74_c1;
  assign nS_st5_b75_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b75_c0 : nS_st4_b75_c1;
  assign nS_st5_b76_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b76_c0 : nS_st4_b76_c1;
  assign nS_st5_b77_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b77_c0 : nS_st4_b77_c1;
  assign nS_st5_b78_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b78_c0 : nS_st4_b78_c1;
  assign nS_st5_b79_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b79_c0 : nS_st4_b79_c1;
  assign nS_st5_b80_c1 = nS_st4_b80_c1;
  assign nS_st5_b81_c1 = nS_st4_b81_c1;
  assign nS_st5_b82_c1 = nS_st4_b82_c1;
  assign nS_st5_b83_c1 = nS_st4_b83_c1;
  assign nS_st5_b84_c1 = nS_st4_b84_c1;
  assign nS_st5_b85_c1 = nS_st4_b85_c1;
  assign nS_st5_b86_c1 = nS_st4_b86_c1;
  assign nS_st5_b87_c1 = nS_st4_b87_c1;
  assign nS_st5_b88_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b88_c0 : nS_st4_b88_c1;
  assign nS_st5_b89_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b89_c0 : nS_st4_b89_c1;
  assign nS_st5_b90_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b90_c0 : nS_st4_b90_c1;
  assign nS_st5_b91_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b91_c0 : nS_st4_b91_c1;
  assign nS_st5_b92_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b92_c0 : nS_st4_b92_c1;
  assign nS_st5_b93_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b93_c0 : nS_st4_b93_c1;
  assign nS_st5_b94_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b94_c0 : nS_st4_b94_c1;
  assign nS_st5_b95_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b95_c0 : nS_st4_b95_c1;
  assign nS_st5_b96_c1 = nS_st4_b96_c1;
  assign nS_st5_b97_c1 = nS_st4_b97_c1;
  assign nS_st5_b98_c1 = nS_st4_b98_c1;
  assign nS_st5_b99_c1 = nS_st4_b99_c1;
  assign nS_st5_b100_c1 = nS_st4_b100_c1;
  assign nS_st5_b101_c1 = nS_st4_b101_c1;
  assign nS_st5_b102_c1 = nS_st4_b102_c1;
  assign nS_st5_b103_c1 = nS_st4_b103_c1;
  assign nS_st5_b104_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b104_c0 : nS_st4_b104_c1;
  assign nS_st5_b105_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b105_c0 : nS_st4_b105_c1;
  assign nS_st5_b106_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b106_c0 : nS_st4_b106_c1;
  assign nS_st5_b107_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b107_c0 : nS_st4_b107_c1;
  assign nS_st5_b108_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b108_c0 : nS_st4_b108_c1;
  assign nS_st5_b109_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b109_c0 : nS_st4_b109_c1;
  assign nS_st5_b110_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b110_c0 : nS_st4_b110_c1;
  assign nS_st5_b111_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b111_c0 : nS_st4_b111_c1;
  assign nS_st5_b112_c1 = nS_st4_b112_c1;
  assign nS_st5_b113_c1 = nS_st4_b113_c1;
  assign nS_st5_b114_c1 = nS_st4_b114_c1;
  assign nS_st5_b115_c1 = nS_st4_b115_c1;
  assign nS_st5_b116_c1 = nS_st4_b116_c1;
  assign nS_st5_b117_c1 = nS_st4_b117_c1;
  assign nS_st5_b118_c1 = nS_st4_b118_c1;
  assign nS_st5_b119_c1 = nS_st4_b119_c1;
  assign nS_st5_b120_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b120_c0 : nS_st4_b120_c1;
  assign nS_st5_b121_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b121_c0 : nS_st4_b121_c1;
  assign nS_st5_b122_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b122_c0 : nS_st4_b122_c1;
  assign nS_st5_b123_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b123_c0 : nS_st4_b123_c1;
  assign nS_st5_b124_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b124_c0 : nS_st4_b124_c1;
  assign nS_st5_b125_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b125_c0 : nS_st4_b125_c1;
  assign nS_st5_b126_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b126_c0 : nS_st4_b126_c1;
  assign nS_st5_b127_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b127_c0 : nS_st4_b127_c1;
  assign nS_st5_b128_c1 = nS_st4_b128_c1;
  assign nS_st5_b129_c1 = nS_st4_b129_c1;
  assign nS_st5_b130_c1 = nS_st4_b130_c1;
  assign nS_st5_b131_c1 = nS_st4_b131_c1;
  assign nS_st5_b132_c1 = nS_st4_b132_c1;
  assign nS_st5_b133_c1 = nS_st4_b133_c1;
  assign nS_st5_b134_c1 = nS_st4_b134_c1;
  assign nS_st5_b135_c1 = nS_st4_b135_c1;
  assign nS_st5_b136_c1 = (nC_st4_b135_c1 == 0) ? nS_st4_b136_c0 : nS_st4_b136_c1;
  assign nS_st5_b137_c1 = (nC_st4_b135_c1 == 0) ? nS_st4_b137_c0 : nS_st4_b137_c1;
  assign nS_st5_b138_c1 = (nC_st4_b135_c1 == 0) ? nS_st4_b138_c0 : nS_st4_b138_c1;
  assign nS_st5_b139_c1 = (nC_st4_b135_c1 == 0) ? nS_st4_b139_c0 : nS_st4_b139_c1;
  assign nS_st5_b140_c1 = (nC_st4_b135_c1 == 0) ? nS_st4_b140_c0 : nS_st4_b140_c1;
  assign nS_st5_b141_c1 = (nC_st4_b135_c1 == 0) ? nS_st4_b141_c0 : nS_st4_b141_c1;
  assign nS_st5_b142_c1 = (nC_st4_b135_c1 == 0) ? nS_st4_b142_c0 : nS_st4_b142_c1;
  assign nS_st5_b143_c1 = (nC_st4_b135_c1 == 0) ? nS_st4_b143_c0 : nS_st4_b143_c1;
  assign nS_st5_b144_c1 = nS_st4_b144_c1;
  assign nS_st5_b145_c1 = nS_st4_b145_c1;
  assign nS_st5_b146_c1 = nS_st4_b146_c1;
  assign nS_st5_b147_c1 = nS_st4_b147_c1;
  assign nS_st5_b148_c1 = nS_st4_b148_c1;
  assign nS_st5_b149_c1 = nS_st4_b149_c1;
  assign nS_st5_b150_c1 = nS_st4_b150_c1;
  assign nS_st5_b151_c1 = nS_st4_b151_c1;
  assign nS_st5_b152_c1 = (nC_st4_b151_c1 == 0) ? nS_st4_b152_c0 : nS_st4_b152_c1;
  assign nS_st5_b153_c1 = (nC_st4_b151_c1 == 0) ? nS_st4_b153_c0 : nS_st4_b153_c1;
  assign nS_st5_b154_c1 = (nC_st4_b151_c1 == 0) ? nS_st4_b154_c0 : nS_st4_b154_c1;
  assign nS_st5_b155_c1 = (nC_st4_b151_c1 == 0) ? nS_st4_b155_c0 : nS_st4_b155_c1;
  assign nS_st5_b156_c1 = (nC_st4_b151_c1 == 0) ? nS_st4_b156_c0 : nS_st4_b156_c1;
  assign nS_st5_b157_c1 = (nC_st4_b151_c1 == 0) ? nS_st4_b157_c0 : nS_st4_b157_c1;
  assign nS_st5_b158_c1 = (nC_st4_b151_c1 == 0) ? nS_st4_b158_c0 : nS_st4_b158_c1;
  assign nS_st5_b159_c1 = (nC_st4_b151_c1 == 0) ? nS_st4_b159_c0 : nS_st4_b159_c1;
  assign nS_st5_b160_c1 = nS_st4_b160_c1;
  assign nS_st5_b161_c1 = nS_st4_b161_c1;
  assign nS_st5_b162_c1 = nS_st4_b162_c1;
  assign nS_st5_b163_c1 = nS_st4_b163_c1;
  assign nS_st5_b164_c1 = nS_st4_b164_c1;
  assign nS_st5_b165_c1 = nS_st4_b165_c1;
  assign nS_st5_b166_c1 = nS_st4_b166_c1;
  assign nS_st5_b167_c1 = nS_st4_b167_c1;
  assign nS_st5_b168_c1 = (nC_st4_b167_c1 == 0) ? nS_st4_b168_c0 : nS_st4_b168_c1;
  assign nS_st5_b169_c1 = (nC_st4_b167_c1 == 0) ? nS_st4_b169_c0 : nS_st4_b169_c1;
  assign nS_st5_b170_c1 = (nC_st4_b167_c1 == 0) ? nS_st4_b170_c0 : nS_st4_b170_c1;
  assign nS_st5_b171_c1 = (nC_st4_b167_c1 == 0) ? nS_st4_b171_c0 : nS_st4_b171_c1;
  assign nS_st5_b172_c1 = (nC_st4_b167_c1 == 0) ? nS_st4_b172_c0 : nS_st4_b172_c1;
  assign nS_st5_b173_c1 = (nC_st4_b167_c1 == 0) ? nS_st4_b173_c0 : nS_st4_b173_c1;
  assign nS_st5_b174_c1 = (nC_st4_b167_c1 == 0) ? nS_st4_b174_c0 : nS_st4_b174_c1;
  assign nS_st5_b175_c1 = (nC_st4_b167_c1 == 0) ? nS_st4_b175_c0 : nS_st4_b175_c1;
  assign nS_st5_b176_c1 = nS_st4_b176_c1;
  assign nS_st5_b177_c1 = nS_st4_b177_c1;
  assign nS_st5_b178_c1 = nS_st4_b178_c1;
  assign nS_st5_b179_c1 = nS_st4_b179_c1;
  assign nS_st5_b180_c1 = nS_st4_b180_c1;
  assign nS_st5_b181_c1 = nS_st4_b181_c1;
  assign nS_st5_b182_c1 = nS_st4_b182_c1;
  assign nS_st5_b183_c1 = nS_st4_b183_c1;
  assign nS_st5_b184_c1 = (nC_st4_b183_c1 == 0) ? nS_st4_b184_c0 : nS_st4_b184_c1;
  assign nS_st5_b185_c1 = (nC_st4_b183_c1 == 0) ? nS_st4_b185_c0 : nS_st4_b185_c1;
  assign nS_st5_b186_c1 = (nC_st4_b183_c1 == 0) ? nS_st4_b186_c0 : nS_st4_b186_c1;
  assign nS_st5_b187_c1 = (nC_st4_b183_c1 == 0) ? nS_st4_b187_c0 : nS_st4_b187_c1;
  assign nS_st5_b188_c1 = (nC_st4_b183_c1 == 0) ? nS_st4_b188_c0 : nS_st4_b188_c1;
  assign nS_st5_b189_c1 = (nC_st4_b183_c1 == 0) ? nS_st4_b189_c0 : nS_st4_b189_c1;
  assign nS_st5_b190_c1 = (nC_st4_b183_c1 == 0) ? nS_st4_b190_c0 : nS_st4_b190_c1;
  assign nS_st5_b191_c1 = (nC_st4_b183_c1 == 0) ? nS_st4_b191_c0 : nS_st4_b191_c1;
  assign nS_st5_b192_c1 = nS_st4_b192_c1;
  assign nS_st5_b193_c1 = nS_st4_b193_c1;
  assign nS_st5_b194_c1 = nS_st4_b194_c1;
  assign nS_st5_b195_c1 = nS_st4_b195_c1;
  assign nS_st5_b196_c1 = nS_st4_b196_c1;
  assign nS_st5_b197_c1 = nS_st4_b197_c1;
  assign nS_st5_b198_c1 = nS_st4_b198_c1;
  assign nS_st5_b199_c1 = nS_st4_b199_c1;
  assign nS_st5_b200_c1 = (nC_st4_b199_c1 == 0) ? nS_st4_b200_c0 : nS_st4_b200_c1;
  assign nS_st5_b201_c1 = (nC_st4_b199_c1 == 0) ? nS_st4_b201_c0 : nS_st4_b201_c1;
  assign nS_st5_b202_c1 = (nC_st4_b199_c1 == 0) ? nS_st4_b202_c0 : nS_st4_b202_c1;
  assign nS_st5_b203_c1 = (nC_st4_b199_c1 == 0) ? nS_st4_b203_c0 : nS_st4_b203_c1;
  assign nS_st5_b204_c1 = (nC_st4_b199_c1 == 0) ? nS_st4_b204_c0 : nS_st4_b204_c1;
  assign nS_st5_b205_c1 = (nC_st4_b199_c1 == 0) ? nS_st4_b205_c0 : nS_st4_b205_c1;
  assign nS_st5_b206_c1 = (nC_st4_b199_c1 == 0) ? nS_st4_b206_c0 : nS_st4_b206_c1;
  assign nS_st5_b207_c1 = (nC_st4_b199_c1 == 0) ? nS_st4_b207_c0 : nS_st4_b207_c1;
  assign nS_st5_b208_c1 = nS_st4_b208_c1;
  assign nS_st5_b209_c1 = nS_st4_b209_c1;
  assign nS_st5_b210_c1 = nS_st4_b210_c1;
  assign nS_st5_b211_c1 = nS_st4_b211_c1;
  assign nS_st5_b212_c1 = nS_st4_b212_c1;
  assign nS_st5_b213_c1 = nS_st4_b213_c1;
  assign nS_st5_b214_c1 = nS_st4_b214_c1;
  assign nS_st5_b215_c1 = nS_st4_b215_c1;
  assign nS_st5_b216_c1 = (nC_st4_b215_c1 == 0) ? nS_st4_b216_c0 : nS_st4_b216_c1;
  assign nS_st5_b217_c1 = (nC_st4_b215_c1 == 0) ? nS_st4_b217_c0 : nS_st4_b217_c1;
  assign nS_st5_b218_c1 = (nC_st4_b215_c1 == 0) ? nS_st4_b218_c0 : nS_st4_b218_c1;
  assign nS_st5_b219_c1 = (nC_st4_b215_c1 == 0) ? nS_st4_b219_c0 : nS_st4_b219_c1;
  assign nS_st5_b220_c1 = (nC_st4_b215_c1 == 0) ? nS_st4_b220_c0 : nS_st4_b220_c1;
  assign nS_st5_b221_c1 = (nC_st4_b215_c1 == 0) ? nS_st4_b221_c0 : nS_st4_b221_c1;
  assign nS_st5_b222_c1 = (nC_st4_b215_c1 == 0) ? nS_st4_b222_c0 : nS_st4_b222_c1;
  assign nS_st5_b223_c1 = (nC_st4_b215_c1 == 0) ? nS_st4_b223_c0 : nS_st4_b223_c1;
  assign nS_st5_b224_c1 = nS_st4_b224_c1;
  assign nS_st5_b225_c1 = nS_st4_b225_c1;
  assign nS_st5_b226_c1 = nS_st4_b226_c1;
  assign nS_st5_b227_c1 = nS_st4_b227_c1;
  assign nS_st5_b228_c1 = nS_st4_b228_c1;
  assign nS_st5_b229_c1 = nS_st4_b229_c1;
  assign nS_st5_b230_c1 = nS_st4_b230_c1;
  assign nS_st5_b231_c1 = nS_st4_b231_c1;
  assign nS_st5_b232_c1 = (nC_st4_b231_c1 == 0) ? nS_st4_b232_c0 : nS_st4_b232_c1;
  assign nS_st5_b233_c1 = (nC_st4_b231_c1 == 0) ? nS_st4_b233_c0 : nS_st4_b233_c1;
  assign nS_st5_b234_c1 = (nC_st4_b231_c1 == 0) ? nS_st4_b234_c0 : nS_st4_b234_c1;
  assign nS_st5_b235_c1 = (nC_st4_b231_c1 == 0) ? nS_st4_b235_c0 : nS_st4_b235_c1;
  assign nS_st5_b236_c1 = (nC_st4_b231_c1 == 0) ? nS_st4_b236_c0 : nS_st4_b236_c1;
  assign nS_st5_b237_c1 = (nC_st4_b231_c1 == 0) ? nS_st4_b237_c0 : nS_st4_b237_c1;
  assign nS_st5_b238_c1 = (nC_st4_b231_c1 == 0) ? nS_st4_b238_c0 : nS_st4_b238_c1;
  assign nS_st5_b239_c1 = (nC_st4_b231_c1 == 0) ? nS_st4_b239_c0 : nS_st4_b239_c1;
  assign nS_st5_b240_c1 = nS_st4_b240_c1;
  assign nS_st5_b241_c1 = nS_st4_b241_c1;
  assign nS_st5_b242_c1 = nS_st4_b242_c1;
  assign nS_st5_b243_c1 = nS_st4_b243_c1;
  assign nS_st5_b244_c1 = nS_st4_b244_c1;
  assign nS_st5_b245_c1 = nS_st4_b245_c1;
  assign nS_st5_b246_c1 = nS_st4_b246_c1;
  assign nS_st5_b247_c1 = nS_st4_b247_c1;
  assign nS_st5_b248_c1 = (nC_st4_b247_c1 == 0) ? nS_st4_b248_c0 : nS_st4_b248_c1;
  assign nS_st5_b249_c1 = (nC_st4_b247_c1 == 0) ? nS_st4_b249_c0 : nS_st4_b249_c1;
  assign nS_st5_b250_c1 = (nC_st4_b247_c1 == 0) ? nS_st4_b250_c0 : nS_st4_b250_c1;
  assign nS_st5_b251_c1 = (nC_st4_b247_c1 == 0) ? nS_st4_b251_c0 : nS_st4_b251_c1;
  assign nS_st5_b252_c1 = (nC_st4_b247_c1 == 0) ? nS_st4_b252_c0 : nS_st4_b252_c1;
  assign nS_st5_b253_c1 = (nC_st4_b247_c1 == 0) ? nS_st4_b253_c0 : nS_st4_b253_c1;
  assign nS_st5_b254_c1 = (nC_st4_b247_c1 == 0) ? nS_st4_b254_c0 : nS_st4_b254_c1;
  assign nS_st5_b255_c1 = (nC_st4_b247_c1 == 0) ? nS_st4_b255_c0 : nS_st4_b255_c1;
  assign nC_st5_b15_c0 = (nC_st4_b7_c0 == 0) ? nC_st4_b15_c0 : nC_st4_b15_c1;
  assign nC_st5_b31_c0 = (nC_st4_b23_c0 == 0) ? nC_st4_b31_c0 : nC_st4_b31_c1;
  assign nC_st5_b47_c0 = (nC_st4_b39_c0 == 0) ? nC_st4_b47_c0 : nC_st4_b47_c1;
  assign nC_st5_b63_c0 = (nC_st4_b55_c0 == 0) ? nC_st4_b63_c0 : nC_st4_b63_c1;
  assign nC_st5_b79_c0 = (nC_st4_b71_c0 == 0) ? nC_st4_b79_c0 : nC_st4_b79_c1;
  assign nC_st5_b95_c0 = (nC_st4_b87_c0 == 0) ? nC_st4_b95_c0 : nC_st4_b95_c1;
  assign nC_st5_b111_c0 = (nC_st4_b103_c0 == 0) ? nC_st4_b111_c0 : nC_st4_b111_c1;
  assign nC_st5_b127_c0 = (nC_st4_b119_c0 == 0) ? nC_st4_b127_c0 : nC_st4_b127_c1;
  assign nC_st5_b143_c0 = (nC_st4_b135_c0 == 0) ? nC_st4_b143_c0 : nC_st4_b143_c1;
  assign nC_st5_b159_c0 = (nC_st4_b151_c0 == 0) ? nC_st4_b159_c0 : nC_st4_b159_c1;
  assign nC_st5_b175_c0 = (nC_st4_b167_c0 == 0) ? nC_st4_b175_c0 : nC_st4_b175_c1;
  assign nC_st5_b191_c0 = (nC_st4_b183_c0 == 0) ? nC_st4_b191_c0 : nC_st4_b191_c1;
  assign nC_st5_b207_c0 = (nC_st4_b199_c0 == 0) ? nC_st4_b207_c0 : nC_st4_b207_c1;
  assign nC_st5_b223_c0 = (nC_st4_b215_c0 == 0) ? nC_st4_b223_c0 : nC_st4_b223_c1;
  assign nC_st5_b239_c0 = (nC_st4_b231_c0 == 0) ? nC_st4_b239_c0 : nC_st4_b239_c1;
  assign nC_st5_b255_c0 = (nC_st4_b247_c0 == 0) ? nC_st4_b255_c0 : nC_st4_b255_c1;
  assign nC_st5_b15_c1 = (nC_st4_b7_c1 == 0) ? nC_st4_b15_c0 : nC_st4_b15_c1;
  assign nC_st5_b31_c1 = (nC_st4_b23_c1 == 0) ? nC_st4_b31_c0 : nC_st4_b31_c1;
  assign nC_st5_b47_c1 = (nC_st4_b39_c1 == 0) ? nC_st4_b47_c0 : nC_st4_b47_c1;
  assign nC_st5_b63_c1 = (nC_st4_b55_c1 == 0) ? nC_st4_b63_c0 : nC_st4_b63_c1;
  assign nC_st5_b79_c1 = (nC_st4_b71_c1 == 0) ? nC_st4_b79_c0 : nC_st4_b79_c1;
  assign nC_st5_b95_c1 = (nC_st4_b87_c1 == 0) ? nC_st4_b95_c0 : nC_st4_b95_c1;
  assign nC_st5_b111_c1 = (nC_st4_b103_c1 == 0) ? nC_st4_b111_c0 : nC_st4_b111_c1;
  assign nC_st5_b127_c1 = (nC_st4_b119_c1 == 0) ? nC_st4_b127_c0 : nC_st4_b127_c1;
  assign nC_st5_b143_c1 = (nC_st4_b135_c1 == 0) ? nC_st4_b143_c0 : nC_st4_b143_c1;
  assign nC_st5_b159_c1 = (nC_st4_b151_c1 == 0) ? nC_st4_b159_c0 : nC_st4_b159_c1;
  assign nC_st5_b175_c1 = (nC_st4_b167_c1 == 0) ? nC_st4_b175_c0 : nC_st4_b175_c1;
  assign nC_st5_b191_c1 = (nC_st4_b183_c1 == 0) ? nC_st4_b191_c0 : nC_st4_b191_c1;
  assign nC_st5_b207_c1 = (nC_st4_b199_c1 == 0) ? nC_st4_b207_c0 : nC_st4_b207_c1;
  assign nC_st5_b223_c1 = (nC_st4_b215_c1 == 0) ? nC_st4_b223_c0 : nC_st4_b223_c1;
  assign nC_st5_b239_c1 = (nC_st4_b231_c1 == 0) ? nC_st4_b239_c0 : nC_st4_b239_c1;
  assign nC_st5_b255_c1 = (nC_st4_b247_c1 == 0) ? nC_st4_b255_c0 : nC_st4_b255_c1;

  assign nS_st6_b0_c0 = nS_st5_b0_c0;
  assign nS_st6_b1_c0 = nS_st5_b1_c0;
  assign nS_st6_b2_c0 = nS_st5_b2_c0;
  assign nS_st6_b3_c0 = nS_st5_b3_c0;
  assign nS_st6_b4_c0 = nS_st5_b4_c0;
  assign nS_st6_b5_c0 = nS_st5_b5_c0;
  assign nS_st6_b6_c0 = nS_st5_b6_c0;
  assign nS_st6_b7_c0 = nS_st5_b7_c0;
  assign nS_st6_b8_c0 = nS_st5_b8_c0;
  assign nS_st6_b9_c0 = nS_st5_b9_c0;
  assign nS_st6_b10_c0 = nS_st5_b10_c0;
  assign nS_st6_b11_c0 = nS_st5_b11_c0;
  assign nS_st6_b12_c0 = nS_st5_b12_c0;
  assign nS_st6_b13_c0 = nS_st5_b13_c0;
  assign nS_st6_b14_c0 = nS_st5_b14_c0;
  assign nS_st6_b15_c0 = nS_st5_b15_c0;
  assign nS_st6_b16_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b16_c0 : nS_st5_b16_c1;
  assign nS_st6_b17_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b17_c0 : nS_st5_b17_c1;
  assign nS_st6_b18_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b18_c0 : nS_st5_b18_c1;
  assign nS_st6_b19_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b19_c0 : nS_st5_b19_c1;
  assign nS_st6_b20_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b20_c0 : nS_st5_b20_c1;
  assign nS_st6_b21_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b21_c0 : nS_st5_b21_c1;
  assign nS_st6_b22_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b22_c0 : nS_st5_b22_c1;
  assign nS_st6_b23_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b23_c0 : nS_st5_b23_c1;
  assign nS_st6_b24_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b24_c0 : nS_st5_b24_c1;
  assign nS_st6_b25_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b25_c0 : nS_st5_b25_c1;
  assign nS_st6_b26_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b26_c0 : nS_st5_b26_c1;
  assign nS_st6_b27_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b27_c0 : nS_st5_b27_c1;
  assign nS_st6_b28_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b28_c0 : nS_st5_b28_c1;
  assign nS_st6_b29_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b29_c0 : nS_st5_b29_c1;
  assign nS_st6_b30_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b30_c0 : nS_st5_b30_c1;
  assign nS_st6_b31_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b31_c0 : nS_st5_b31_c1;
  assign nS_st6_b32_c0 = nS_st5_b32_c0;
  assign nS_st6_b33_c0 = nS_st5_b33_c0;
  assign nS_st6_b34_c0 = nS_st5_b34_c0;
  assign nS_st6_b35_c0 = nS_st5_b35_c0;
  assign nS_st6_b36_c0 = nS_st5_b36_c0;
  assign nS_st6_b37_c0 = nS_st5_b37_c0;
  assign nS_st6_b38_c0 = nS_st5_b38_c0;
  assign nS_st6_b39_c0 = nS_st5_b39_c0;
  assign nS_st6_b40_c0 = nS_st5_b40_c0;
  assign nS_st6_b41_c0 = nS_st5_b41_c0;
  assign nS_st6_b42_c0 = nS_st5_b42_c0;
  assign nS_st6_b43_c0 = nS_st5_b43_c0;
  assign nS_st6_b44_c0 = nS_st5_b44_c0;
  assign nS_st6_b45_c0 = nS_st5_b45_c0;
  assign nS_st6_b46_c0 = nS_st5_b46_c0;
  assign nS_st6_b47_c0 = nS_st5_b47_c0;
  assign nS_st6_b48_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b48_c0 : nS_st5_b48_c1;
  assign nS_st6_b49_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b49_c0 : nS_st5_b49_c1;
  assign nS_st6_b50_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b50_c0 : nS_st5_b50_c1;
  assign nS_st6_b51_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b51_c0 : nS_st5_b51_c1;
  assign nS_st6_b52_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b52_c0 : nS_st5_b52_c1;
  assign nS_st6_b53_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b53_c0 : nS_st5_b53_c1;
  assign nS_st6_b54_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b54_c0 : nS_st5_b54_c1;
  assign nS_st6_b55_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b55_c0 : nS_st5_b55_c1;
  assign nS_st6_b56_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b56_c0 : nS_st5_b56_c1;
  assign nS_st6_b57_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b57_c0 : nS_st5_b57_c1;
  assign nS_st6_b58_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b58_c0 : nS_st5_b58_c1;
  assign nS_st6_b59_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b59_c0 : nS_st5_b59_c1;
  assign nS_st6_b60_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b60_c0 : nS_st5_b60_c1;
  assign nS_st6_b61_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b61_c0 : nS_st5_b61_c1;
  assign nS_st6_b62_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b62_c0 : nS_st5_b62_c1;
  assign nS_st6_b63_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b63_c0 : nS_st5_b63_c1;
  assign nS_st6_b64_c0 = nS_st5_b64_c0;
  assign nS_st6_b65_c0 = nS_st5_b65_c0;
  assign nS_st6_b66_c0 = nS_st5_b66_c0;
  assign nS_st6_b67_c0 = nS_st5_b67_c0;
  assign nS_st6_b68_c0 = nS_st5_b68_c0;
  assign nS_st6_b69_c0 = nS_st5_b69_c0;
  assign nS_st6_b70_c0 = nS_st5_b70_c0;
  assign nS_st6_b71_c0 = nS_st5_b71_c0;
  assign nS_st6_b72_c0 = nS_st5_b72_c0;
  assign nS_st6_b73_c0 = nS_st5_b73_c0;
  assign nS_st6_b74_c0 = nS_st5_b74_c0;
  assign nS_st6_b75_c0 = nS_st5_b75_c0;
  assign nS_st6_b76_c0 = nS_st5_b76_c0;
  assign nS_st6_b77_c0 = nS_st5_b77_c0;
  assign nS_st6_b78_c0 = nS_st5_b78_c0;
  assign nS_st6_b79_c0 = nS_st5_b79_c0;
  assign nS_st6_b80_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b80_c0 : nS_st5_b80_c1;
  assign nS_st6_b81_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b81_c0 : nS_st5_b81_c1;
  assign nS_st6_b82_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b82_c0 : nS_st5_b82_c1;
  assign nS_st6_b83_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b83_c0 : nS_st5_b83_c1;
  assign nS_st6_b84_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b84_c0 : nS_st5_b84_c1;
  assign nS_st6_b85_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b85_c0 : nS_st5_b85_c1;
  assign nS_st6_b86_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b86_c0 : nS_st5_b86_c1;
  assign nS_st6_b87_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b87_c0 : nS_st5_b87_c1;
  assign nS_st6_b88_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b88_c0 : nS_st5_b88_c1;
  assign nS_st6_b89_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b89_c0 : nS_st5_b89_c1;
  assign nS_st6_b90_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b90_c0 : nS_st5_b90_c1;
  assign nS_st6_b91_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b91_c0 : nS_st5_b91_c1;
  assign nS_st6_b92_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b92_c0 : nS_st5_b92_c1;
  assign nS_st6_b93_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b93_c0 : nS_st5_b93_c1;
  assign nS_st6_b94_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b94_c0 : nS_st5_b94_c1;
  assign nS_st6_b95_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b95_c0 : nS_st5_b95_c1;
  assign nS_st6_b96_c0 = nS_st5_b96_c0;
  assign nS_st6_b97_c0 = nS_st5_b97_c0;
  assign nS_st6_b98_c0 = nS_st5_b98_c0;
  assign nS_st6_b99_c0 = nS_st5_b99_c0;
  assign nS_st6_b100_c0 = nS_st5_b100_c0;
  assign nS_st6_b101_c0 = nS_st5_b101_c0;
  assign nS_st6_b102_c0 = nS_st5_b102_c0;
  assign nS_st6_b103_c0 = nS_st5_b103_c0;
  assign nS_st6_b104_c0 = nS_st5_b104_c0;
  assign nS_st6_b105_c0 = nS_st5_b105_c0;
  assign nS_st6_b106_c0 = nS_st5_b106_c0;
  assign nS_st6_b107_c0 = nS_st5_b107_c0;
  assign nS_st6_b108_c0 = nS_st5_b108_c0;
  assign nS_st6_b109_c0 = nS_st5_b109_c0;
  assign nS_st6_b110_c0 = nS_st5_b110_c0;
  assign nS_st6_b111_c0 = nS_st5_b111_c0;
  assign nS_st6_b112_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b112_c0 : nS_st5_b112_c1;
  assign nS_st6_b113_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b113_c0 : nS_st5_b113_c1;
  assign nS_st6_b114_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b114_c0 : nS_st5_b114_c1;
  assign nS_st6_b115_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b115_c0 : nS_st5_b115_c1;
  assign nS_st6_b116_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b116_c0 : nS_st5_b116_c1;
  assign nS_st6_b117_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b117_c0 : nS_st5_b117_c1;
  assign nS_st6_b118_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b118_c0 : nS_st5_b118_c1;
  assign nS_st6_b119_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b119_c0 : nS_st5_b119_c1;
  assign nS_st6_b120_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b120_c0 : nS_st5_b120_c1;
  assign nS_st6_b121_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b121_c0 : nS_st5_b121_c1;
  assign nS_st6_b122_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b122_c0 : nS_st5_b122_c1;
  assign nS_st6_b123_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b123_c0 : nS_st5_b123_c1;
  assign nS_st6_b124_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b124_c0 : nS_st5_b124_c1;
  assign nS_st6_b125_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b125_c0 : nS_st5_b125_c1;
  assign nS_st6_b126_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b126_c0 : nS_st5_b126_c1;
  assign nS_st6_b127_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b127_c0 : nS_st5_b127_c1;
  assign nS_st6_b128_c0 = nS_st5_b128_c0;
  assign nS_st6_b129_c0 = nS_st5_b129_c0;
  assign nS_st6_b130_c0 = nS_st5_b130_c0;
  assign nS_st6_b131_c0 = nS_st5_b131_c0;
  assign nS_st6_b132_c0 = nS_st5_b132_c0;
  assign nS_st6_b133_c0 = nS_st5_b133_c0;
  assign nS_st6_b134_c0 = nS_st5_b134_c0;
  assign nS_st6_b135_c0 = nS_st5_b135_c0;
  assign nS_st6_b136_c0 = nS_st5_b136_c0;
  assign nS_st6_b137_c0 = nS_st5_b137_c0;
  assign nS_st6_b138_c0 = nS_st5_b138_c0;
  assign nS_st6_b139_c0 = nS_st5_b139_c0;
  assign nS_st6_b140_c0 = nS_st5_b140_c0;
  assign nS_st6_b141_c0 = nS_st5_b141_c0;
  assign nS_st6_b142_c0 = nS_st5_b142_c0;
  assign nS_st6_b143_c0 = nS_st5_b143_c0;
  assign nS_st6_b144_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b144_c0 : nS_st5_b144_c1;
  assign nS_st6_b145_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b145_c0 : nS_st5_b145_c1;
  assign nS_st6_b146_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b146_c0 : nS_st5_b146_c1;
  assign nS_st6_b147_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b147_c0 : nS_st5_b147_c1;
  assign nS_st6_b148_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b148_c0 : nS_st5_b148_c1;
  assign nS_st6_b149_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b149_c0 : nS_st5_b149_c1;
  assign nS_st6_b150_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b150_c0 : nS_st5_b150_c1;
  assign nS_st6_b151_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b151_c0 : nS_st5_b151_c1;
  assign nS_st6_b152_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b152_c0 : nS_st5_b152_c1;
  assign nS_st6_b153_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b153_c0 : nS_st5_b153_c1;
  assign nS_st6_b154_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b154_c0 : nS_st5_b154_c1;
  assign nS_st6_b155_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b155_c0 : nS_st5_b155_c1;
  assign nS_st6_b156_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b156_c0 : nS_st5_b156_c1;
  assign nS_st6_b157_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b157_c0 : nS_st5_b157_c1;
  assign nS_st6_b158_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b158_c0 : nS_st5_b158_c1;
  assign nS_st6_b159_c0 = (nC_st5_b143_c0 == 0) ? nS_st5_b159_c0 : nS_st5_b159_c1;
  assign nS_st6_b160_c0 = nS_st5_b160_c0;
  assign nS_st6_b161_c0 = nS_st5_b161_c0;
  assign nS_st6_b162_c0 = nS_st5_b162_c0;
  assign nS_st6_b163_c0 = nS_st5_b163_c0;
  assign nS_st6_b164_c0 = nS_st5_b164_c0;
  assign nS_st6_b165_c0 = nS_st5_b165_c0;
  assign nS_st6_b166_c0 = nS_st5_b166_c0;
  assign nS_st6_b167_c0 = nS_st5_b167_c0;
  assign nS_st6_b168_c0 = nS_st5_b168_c0;
  assign nS_st6_b169_c0 = nS_st5_b169_c0;
  assign nS_st6_b170_c0 = nS_st5_b170_c0;
  assign nS_st6_b171_c0 = nS_st5_b171_c0;
  assign nS_st6_b172_c0 = nS_st5_b172_c0;
  assign nS_st6_b173_c0 = nS_st5_b173_c0;
  assign nS_st6_b174_c0 = nS_st5_b174_c0;
  assign nS_st6_b175_c0 = nS_st5_b175_c0;
  assign nS_st6_b176_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b176_c0 : nS_st5_b176_c1;
  assign nS_st6_b177_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b177_c0 : nS_st5_b177_c1;
  assign nS_st6_b178_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b178_c0 : nS_st5_b178_c1;
  assign nS_st6_b179_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b179_c0 : nS_st5_b179_c1;
  assign nS_st6_b180_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b180_c0 : nS_st5_b180_c1;
  assign nS_st6_b181_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b181_c0 : nS_st5_b181_c1;
  assign nS_st6_b182_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b182_c0 : nS_st5_b182_c1;
  assign nS_st6_b183_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b183_c0 : nS_st5_b183_c1;
  assign nS_st6_b184_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b184_c0 : nS_st5_b184_c1;
  assign nS_st6_b185_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b185_c0 : nS_st5_b185_c1;
  assign nS_st6_b186_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b186_c0 : nS_st5_b186_c1;
  assign nS_st6_b187_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b187_c0 : nS_st5_b187_c1;
  assign nS_st6_b188_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b188_c0 : nS_st5_b188_c1;
  assign nS_st6_b189_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b189_c0 : nS_st5_b189_c1;
  assign nS_st6_b190_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b190_c0 : nS_st5_b190_c1;
  assign nS_st6_b191_c0 = (nC_st5_b175_c0 == 0) ? nS_st5_b191_c0 : nS_st5_b191_c1;
  assign nS_st6_b192_c0 = nS_st5_b192_c0;
  assign nS_st6_b193_c0 = nS_st5_b193_c0;
  assign nS_st6_b194_c0 = nS_st5_b194_c0;
  assign nS_st6_b195_c0 = nS_st5_b195_c0;
  assign nS_st6_b196_c0 = nS_st5_b196_c0;
  assign nS_st6_b197_c0 = nS_st5_b197_c0;
  assign nS_st6_b198_c0 = nS_st5_b198_c0;
  assign nS_st6_b199_c0 = nS_st5_b199_c0;
  assign nS_st6_b200_c0 = nS_st5_b200_c0;
  assign nS_st6_b201_c0 = nS_st5_b201_c0;
  assign nS_st6_b202_c0 = nS_st5_b202_c0;
  assign nS_st6_b203_c0 = nS_st5_b203_c0;
  assign nS_st6_b204_c0 = nS_st5_b204_c0;
  assign nS_st6_b205_c0 = nS_st5_b205_c0;
  assign nS_st6_b206_c0 = nS_st5_b206_c0;
  assign nS_st6_b207_c0 = nS_st5_b207_c0;
  assign nS_st6_b208_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b208_c0 : nS_st5_b208_c1;
  assign nS_st6_b209_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b209_c0 : nS_st5_b209_c1;
  assign nS_st6_b210_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b210_c0 : nS_st5_b210_c1;
  assign nS_st6_b211_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b211_c0 : nS_st5_b211_c1;
  assign nS_st6_b212_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b212_c0 : nS_st5_b212_c1;
  assign nS_st6_b213_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b213_c0 : nS_st5_b213_c1;
  assign nS_st6_b214_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b214_c0 : nS_st5_b214_c1;
  assign nS_st6_b215_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b215_c0 : nS_st5_b215_c1;
  assign nS_st6_b216_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b216_c0 : nS_st5_b216_c1;
  assign nS_st6_b217_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b217_c0 : nS_st5_b217_c1;
  assign nS_st6_b218_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b218_c0 : nS_st5_b218_c1;
  assign nS_st6_b219_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b219_c0 : nS_st5_b219_c1;
  assign nS_st6_b220_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b220_c0 : nS_st5_b220_c1;
  assign nS_st6_b221_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b221_c0 : nS_st5_b221_c1;
  assign nS_st6_b222_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b222_c0 : nS_st5_b222_c1;
  assign nS_st6_b223_c0 = (nC_st5_b207_c0 == 0) ? nS_st5_b223_c0 : nS_st5_b223_c1;
  assign nS_st6_b224_c0 = nS_st5_b224_c0;
  assign nS_st6_b225_c0 = nS_st5_b225_c0;
  assign nS_st6_b226_c0 = nS_st5_b226_c0;
  assign nS_st6_b227_c0 = nS_st5_b227_c0;
  assign nS_st6_b228_c0 = nS_st5_b228_c0;
  assign nS_st6_b229_c0 = nS_st5_b229_c0;
  assign nS_st6_b230_c0 = nS_st5_b230_c0;
  assign nS_st6_b231_c0 = nS_st5_b231_c0;
  assign nS_st6_b232_c0 = nS_st5_b232_c0;
  assign nS_st6_b233_c0 = nS_st5_b233_c0;
  assign nS_st6_b234_c0 = nS_st5_b234_c0;
  assign nS_st6_b235_c0 = nS_st5_b235_c0;
  assign nS_st6_b236_c0 = nS_st5_b236_c0;
  assign nS_st6_b237_c0 = nS_st5_b237_c0;
  assign nS_st6_b238_c0 = nS_st5_b238_c0;
  assign nS_st6_b239_c0 = nS_st5_b239_c0;
  assign nS_st6_b240_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b240_c0 : nS_st5_b240_c1;
  assign nS_st6_b241_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b241_c0 : nS_st5_b241_c1;
  assign nS_st6_b242_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b242_c0 : nS_st5_b242_c1;
  assign nS_st6_b243_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b243_c0 : nS_st5_b243_c1;
  assign nS_st6_b244_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b244_c0 : nS_st5_b244_c1;
  assign nS_st6_b245_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b245_c0 : nS_st5_b245_c1;
  assign nS_st6_b246_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b246_c0 : nS_st5_b246_c1;
  assign nS_st6_b247_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b247_c0 : nS_st5_b247_c1;
  assign nS_st6_b248_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b248_c0 : nS_st5_b248_c1;
  assign nS_st6_b249_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b249_c0 : nS_st5_b249_c1;
  assign nS_st6_b250_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b250_c0 : nS_st5_b250_c1;
  assign nS_st6_b251_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b251_c0 : nS_st5_b251_c1;
  assign nS_st6_b252_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b252_c0 : nS_st5_b252_c1;
  assign nS_st6_b253_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b253_c0 : nS_st5_b253_c1;
  assign nS_st6_b254_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b254_c0 : nS_st5_b254_c1;
  assign nS_st6_b255_c0 = (nC_st5_b239_c0 == 0) ? nS_st5_b255_c0 : nS_st5_b255_c1;
  assign nS_st6_b0_c1 = nS_st5_b0_c1;
  assign nS_st6_b1_c1 = nS_st5_b1_c1;
  assign nS_st6_b2_c1 = nS_st5_b2_c1;
  assign nS_st6_b3_c1 = nS_st5_b3_c1;
  assign nS_st6_b4_c1 = nS_st5_b4_c1;
  assign nS_st6_b5_c1 = nS_st5_b5_c1;
  assign nS_st6_b6_c1 = nS_st5_b6_c1;
  assign nS_st6_b7_c1 = nS_st5_b7_c1;
  assign nS_st6_b8_c1 = nS_st5_b8_c1;
  assign nS_st6_b9_c1 = nS_st5_b9_c1;
  assign nS_st6_b10_c1 = nS_st5_b10_c1;
  assign nS_st6_b11_c1 = nS_st5_b11_c1;
  assign nS_st6_b12_c1 = nS_st5_b12_c1;
  assign nS_st6_b13_c1 = nS_st5_b13_c1;
  assign nS_st6_b14_c1 = nS_st5_b14_c1;
  assign nS_st6_b15_c1 = nS_st5_b15_c1;
  assign nS_st6_b16_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b16_c0 : nS_st5_b16_c1;
  assign nS_st6_b17_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b17_c0 : nS_st5_b17_c1;
  assign nS_st6_b18_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b18_c0 : nS_st5_b18_c1;
  assign nS_st6_b19_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b19_c0 : nS_st5_b19_c1;
  assign nS_st6_b20_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b20_c0 : nS_st5_b20_c1;
  assign nS_st6_b21_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b21_c0 : nS_st5_b21_c1;
  assign nS_st6_b22_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b22_c0 : nS_st5_b22_c1;
  assign nS_st6_b23_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b23_c0 : nS_st5_b23_c1;
  assign nS_st6_b24_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b24_c0 : nS_st5_b24_c1;
  assign nS_st6_b25_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b25_c0 : nS_st5_b25_c1;
  assign nS_st6_b26_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b26_c0 : nS_st5_b26_c1;
  assign nS_st6_b27_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b27_c0 : nS_st5_b27_c1;
  assign nS_st6_b28_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b28_c0 : nS_st5_b28_c1;
  assign nS_st6_b29_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b29_c0 : nS_st5_b29_c1;
  assign nS_st6_b30_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b30_c0 : nS_st5_b30_c1;
  assign nS_st6_b31_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b31_c0 : nS_st5_b31_c1;
  assign nS_st6_b32_c1 = nS_st5_b32_c1;
  assign nS_st6_b33_c1 = nS_st5_b33_c1;
  assign nS_st6_b34_c1 = nS_st5_b34_c1;
  assign nS_st6_b35_c1 = nS_st5_b35_c1;
  assign nS_st6_b36_c1 = nS_st5_b36_c1;
  assign nS_st6_b37_c1 = nS_st5_b37_c1;
  assign nS_st6_b38_c1 = nS_st5_b38_c1;
  assign nS_st6_b39_c1 = nS_st5_b39_c1;
  assign nS_st6_b40_c1 = nS_st5_b40_c1;
  assign nS_st6_b41_c1 = nS_st5_b41_c1;
  assign nS_st6_b42_c1 = nS_st5_b42_c1;
  assign nS_st6_b43_c1 = nS_st5_b43_c1;
  assign nS_st6_b44_c1 = nS_st5_b44_c1;
  assign nS_st6_b45_c1 = nS_st5_b45_c1;
  assign nS_st6_b46_c1 = nS_st5_b46_c1;
  assign nS_st6_b47_c1 = nS_st5_b47_c1;
  assign nS_st6_b48_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b48_c0 : nS_st5_b48_c1;
  assign nS_st6_b49_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b49_c0 : nS_st5_b49_c1;
  assign nS_st6_b50_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b50_c0 : nS_st5_b50_c1;
  assign nS_st6_b51_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b51_c0 : nS_st5_b51_c1;
  assign nS_st6_b52_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b52_c0 : nS_st5_b52_c1;
  assign nS_st6_b53_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b53_c0 : nS_st5_b53_c1;
  assign nS_st6_b54_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b54_c0 : nS_st5_b54_c1;
  assign nS_st6_b55_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b55_c0 : nS_st5_b55_c1;
  assign nS_st6_b56_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b56_c0 : nS_st5_b56_c1;
  assign nS_st6_b57_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b57_c0 : nS_st5_b57_c1;
  assign nS_st6_b58_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b58_c0 : nS_st5_b58_c1;
  assign nS_st6_b59_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b59_c0 : nS_st5_b59_c1;
  assign nS_st6_b60_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b60_c0 : nS_st5_b60_c1;
  assign nS_st6_b61_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b61_c0 : nS_st5_b61_c1;
  assign nS_st6_b62_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b62_c0 : nS_st5_b62_c1;
  assign nS_st6_b63_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b63_c0 : nS_st5_b63_c1;
  assign nS_st6_b64_c1 = nS_st5_b64_c1;
  assign nS_st6_b65_c1 = nS_st5_b65_c1;
  assign nS_st6_b66_c1 = nS_st5_b66_c1;
  assign nS_st6_b67_c1 = nS_st5_b67_c1;
  assign nS_st6_b68_c1 = nS_st5_b68_c1;
  assign nS_st6_b69_c1 = nS_st5_b69_c1;
  assign nS_st6_b70_c1 = nS_st5_b70_c1;
  assign nS_st6_b71_c1 = nS_st5_b71_c1;
  assign nS_st6_b72_c1 = nS_st5_b72_c1;
  assign nS_st6_b73_c1 = nS_st5_b73_c1;
  assign nS_st6_b74_c1 = nS_st5_b74_c1;
  assign nS_st6_b75_c1 = nS_st5_b75_c1;
  assign nS_st6_b76_c1 = nS_st5_b76_c1;
  assign nS_st6_b77_c1 = nS_st5_b77_c1;
  assign nS_st6_b78_c1 = nS_st5_b78_c1;
  assign nS_st6_b79_c1 = nS_st5_b79_c1;
  assign nS_st6_b80_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b80_c0 : nS_st5_b80_c1;
  assign nS_st6_b81_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b81_c0 : nS_st5_b81_c1;
  assign nS_st6_b82_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b82_c0 : nS_st5_b82_c1;
  assign nS_st6_b83_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b83_c0 : nS_st5_b83_c1;
  assign nS_st6_b84_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b84_c0 : nS_st5_b84_c1;
  assign nS_st6_b85_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b85_c0 : nS_st5_b85_c1;
  assign nS_st6_b86_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b86_c0 : nS_st5_b86_c1;
  assign nS_st6_b87_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b87_c0 : nS_st5_b87_c1;
  assign nS_st6_b88_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b88_c0 : nS_st5_b88_c1;
  assign nS_st6_b89_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b89_c0 : nS_st5_b89_c1;
  assign nS_st6_b90_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b90_c0 : nS_st5_b90_c1;
  assign nS_st6_b91_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b91_c0 : nS_st5_b91_c1;
  assign nS_st6_b92_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b92_c0 : nS_st5_b92_c1;
  assign nS_st6_b93_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b93_c0 : nS_st5_b93_c1;
  assign nS_st6_b94_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b94_c0 : nS_st5_b94_c1;
  assign nS_st6_b95_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b95_c0 : nS_st5_b95_c1;
  assign nS_st6_b96_c1 = nS_st5_b96_c1;
  assign nS_st6_b97_c1 = nS_st5_b97_c1;
  assign nS_st6_b98_c1 = nS_st5_b98_c1;
  assign nS_st6_b99_c1 = nS_st5_b99_c1;
  assign nS_st6_b100_c1 = nS_st5_b100_c1;
  assign nS_st6_b101_c1 = nS_st5_b101_c1;
  assign nS_st6_b102_c1 = nS_st5_b102_c1;
  assign nS_st6_b103_c1 = nS_st5_b103_c1;
  assign nS_st6_b104_c1 = nS_st5_b104_c1;
  assign nS_st6_b105_c1 = nS_st5_b105_c1;
  assign nS_st6_b106_c1 = nS_st5_b106_c1;
  assign nS_st6_b107_c1 = nS_st5_b107_c1;
  assign nS_st6_b108_c1 = nS_st5_b108_c1;
  assign nS_st6_b109_c1 = nS_st5_b109_c1;
  assign nS_st6_b110_c1 = nS_st5_b110_c1;
  assign nS_st6_b111_c1 = nS_st5_b111_c1;
  assign nS_st6_b112_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b112_c0 : nS_st5_b112_c1;
  assign nS_st6_b113_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b113_c0 : nS_st5_b113_c1;
  assign nS_st6_b114_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b114_c0 : nS_st5_b114_c1;
  assign nS_st6_b115_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b115_c0 : nS_st5_b115_c1;
  assign nS_st6_b116_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b116_c0 : nS_st5_b116_c1;
  assign nS_st6_b117_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b117_c0 : nS_st5_b117_c1;
  assign nS_st6_b118_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b118_c0 : nS_st5_b118_c1;
  assign nS_st6_b119_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b119_c0 : nS_st5_b119_c1;
  assign nS_st6_b120_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b120_c0 : nS_st5_b120_c1;
  assign nS_st6_b121_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b121_c0 : nS_st5_b121_c1;
  assign nS_st6_b122_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b122_c0 : nS_st5_b122_c1;
  assign nS_st6_b123_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b123_c0 : nS_st5_b123_c1;
  assign nS_st6_b124_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b124_c0 : nS_st5_b124_c1;
  assign nS_st6_b125_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b125_c0 : nS_st5_b125_c1;
  assign nS_st6_b126_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b126_c0 : nS_st5_b126_c1;
  assign nS_st6_b127_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b127_c0 : nS_st5_b127_c1;
  assign nS_st6_b128_c1 = nS_st5_b128_c1;
  assign nS_st6_b129_c1 = nS_st5_b129_c1;
  assign nS_st6_b130_c1 = nS_st5_b130_c1;
  assign nS_st6_b131_c1 = nS_st5_b131_c1;
  assign nS_st6_b132_c1 = nS_st5_b132_c1;
  assign nS_st6_b133_c1 = nS_st5_b133_c1;
  assign nS_st6_b134_c1 = nS_st5_b134_c1;
  assign nS_st6_b135_c1 = nS_st5_b135_c1;
  assign nS_st6_b136_c1 = nS_st5_b136_c1;
  assign nS_st6_b137_c1 = nS_st5_b137_c1;
  assign nS_st6_b138_c1 = nS_st5_b138_c1;
  assign nS_st6_b139_c1 = nS_st5_b139_c1;
  assign nS_st6_b140_c1 = nS_st5_b140_c1;
  assign nS_st6_b141_c1 = nS_st5_b141_c1;
  assign nS_st6_b142_c1 = nS_st5_b142_c1;
  assign nS_st6_b143_c1 = nS_st5_b143_c1;
  assign nS_st6_b144_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b144_c0 : nS_st5_b144_c1;
  assign nS_st6_b145_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b145_c0 : nS_st5_b145_c1;
  assign nS_st6_b146_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b146_c0 : nS_st5_b146_c1;
  assign nS_st6_b147_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b147_c0 : nS_st5_b147_c1;
  assign nS_st6_b148_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b148_c0 : nS_st5_b148_c1;
  assign nS_st6_b149_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b149_c0 : nS_st5_b149_c1;
  assign nS_st6_b150_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b150_c0 : nS_st5_b150_c1;
  assign nS_st6_b151_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b151_c0 : nS_st5_b151_c1;
  assign nS_st6_b152_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b152_c0 : nS_st5_b152_c1;
  assign nS_st6_b153_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b153_c0 : nS_st5_b153_c1;
  assign nS_st6_b154_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b154_c0 : nS_st5_b154_c1;
  assign nS_st6_b155_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b155_c0 : nS_st5_b155_c1;
  assign nS_st6_b156_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b156_c0 : nS_st5_b156_c1;
  assign nS_st6_b157_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b157_c0 : nS_st5_b157_c1;
  assign nS_st6_b158_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b158_c0 : nS_st5_b158_c1;
  assign nS_st6_b159_c1 = (nC_st5_b143_c1 == 0) ? nS_st5_b159_c0 : nS_st5_b159_c1;
  assign nS_st6_b160_c1 = nS_st5_b160_c1;
  assign nS_st6_b161_c1 = nS_st5_b161_c1;
  assign nS_st6_b162_c1 = nS_st5_b162_c1;
  assign nS_st6_b163_c1 = nS_st5_b163_c1;
  assign nS_st6_b164_c1 = nS_st5_b164_c1;
  assign nS_st6_b165_c1 = nS_st5_b165_c1;
  assign nS_st6_b166_c1 = nS_st5_b166_c1;
  assign nS_st6_b167_c1 = nS_st5_b167_c1;
  assign nS_st6_b168_c1 = nS_st5_b168_c1;
  assign nS_st6_b169_c1 = nS_st5_b169_c1;
  assign nS_st6_b170_c1 = nS_st5_b170_c1;
  assign nS_st6_b171_c1 = nS_st5_b171_c1;
  assign nS_st6_b172_c1 = nS_st5_b172_c1;
  assign nS_st6_b173_c1 = nS_st5_b173_c1;
  assign nS_st6_b174_c1 = nS_st5_b174_c1;
  assign nS_st6_b175_c1 = nS_st5_b175_c1;
  assign nS_st6_b176_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b176_c0 : nS_st5_b176_c1;
  assign nS_st6_b177_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b177_c0 : nS_st5_b177_c1;
  assign nS_st6_b178_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b178_c0 : nS_st5_b178_c1;
  assign nS_st6_b179_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b179_c0 : nS_st5_b179_c1;
  assign nS_st6_b180_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b180_c0 : nS_st5_b180_c1;
  assign nS_st6_b181_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b181_c0 : nS_st5_b181_c1;
  assign nS_st6_b182_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b182_c0 : nS_st5_b182_c1;
  assign nS_st6_b183_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b183_c0 : nS_st5_b183_c1;
  assign nS_st6_b184_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b184_c0 : nS_st5_b184_c1;
  assign nS_st6_b185_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b185_c0 : nS_st5_b185_c1;
  assign nS_st6_b186_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b186_c0 : nS_st5_b186_c1;
  assign nS_st6_b187_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b187_c0 : nS_st5_b187_c1;
  assign nS_st6_b188_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b188_c0 : nS_st5_b188_c1;
  assign nS_st6_b189_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b189_c0 : nS_st5_b189_c1;
  assign nS_st6_b190_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b190_c0 : nS_st5_b190_c1;
  assign nS_st6_b191_c1 = (nC_st5_b175_c1 == 0) ? nS_st5_b191_c0 : nS_st5_b191_c1;
  assign nS_st6_b192_c1 = nS_st5_b192_c1;
  assign nS_st6_b193_c1 = nS_st5_b193_c1;
  assign nS_st6_b194_c1 = nS_st5_b194_c1;
  assign nS_st6_b195_c1 = nS_st5_b195_c1;
  assign nS_st6_b196_c1 = nS_st5_b196_c1;
  assign nS_st6_b197_c1 = nS_st5_b197_c1;
  assign nS_st6_b198_c1 = nS_st5_b198_c1;
  assign nS_st6_b199_c1 = nS_st5_b199_c1;
  assign nS_st6_b200_c1 = nS_st5_b200_c1;
  assign nS_st6_b201_c1 = nS_st5_b201_c1;
  assign nS_st6_b202_c1 = nS_st5_b202_c1;
  assign nS_st6_b203_c1 = nS_st5_b203_c1;
  assign nS_st6_b204_c1 = nS_st5_b204_c1;
  assign nS_st6_b205_c1 = nS_st5_b205_c1;
  assign nS_st6_b206_c1 = nS_st5_b206_c1;
  assign nS_st6_b207_c1 = nS_st5_b207_c1;
  assign nS_st6_b208_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b208_c0 : nS_st5_b208_c1;
  assign nS_st6_b209_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b209_c0 : nS_st5_b209_c1;
  assign nS_st6_b210_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b210_c0 : nS_st5_b210_c1;
  assign nS_st6_b211_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b211_c0 : nS_st5_b211_c1;
  assign nS_st6_b212_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b212_c0 : nS_st5_b212_c1;
  assign nS_st6_b213_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b213_c0 : nS_st5_b213_c1;
  assign nS_st6_b214_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b214_c0 : nS_st5_b214_c1;
  assign nS_st6_b215_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b215_c0 : nS_st5_b215_c1;
  assign nS_st6_b216_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b216_c0 : nS_st5_b216_c1;
  assign nS_st6_b217_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b217_c0 : nS_st5_b217_c1;
  assign nS_st6_b218_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b218_c0 : nS_st5_b218_c1;
  assign nS_st6_b219_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b219_c0 : nS_st5_b219_c1;
  assign nS_st6_b220_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b220_c0 : nS_st5_b220_c1;
  assign nS_st6_b221_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b221_c0 : nS_st5_b221_c1;
  assign nS_st6_b222_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b222_c0 : nS_st5_b222_c1;
  assign nS_st6_b223_c1 = (nC_st5_b207_c1 == 0) ? nS_st5_b223_c0 : nS_st5_b223_c1;
  assign nS_st6_b224_c1 = nS_st5_b224_c1;
  assign nS_st6_b225_c1 = nS_st5_b225_c1;
  assign nS_st6_b226_c1 = nS_st5_b226_c1;
  assign nS_st6_b227_c1 = nS_st5_b227_c1;
  assign nS_st6_b228_c1 = nS_st5_b228_c1;
  assign nS_st6_b229_c1 = nS_st5_b229_c1;
  assign nS_st6_b230_c1 = nS_st5_b230_c1;
  assign nS_st6_b231_c1 = nS_st5_b231_c1;
  assign nS_st6_b232_c1 = nS_st5_b232_c1;
  assign nS_st6_b233_c1 = nS_st5_b233_c1;
  assign nS_st6_b234_c1 = nS_st5_b234_c1;
  assign nS_st6_b235_c1 = nS_st5_b235_c1;
  assign nS_st6_b236_c1 = nS_st5_b236_c1;
  assign nS_st6_b237_c1 = nS_st5_b237_c1;
  assign nS_st6_b238_c1 = nS_st5_b238_c1;
  assign nS_st6_b239_c1 = nS_st5_b239_c1;
  assign nS_st6_b240_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b240_c0 : nS_st5_b240_c1;
  assign nS_st6_b241_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b241_c0 : nS_st5_b241_c1;
  assign nS_st6_b242_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b242_c0 : nS_st5_b242_c1;
  assign nS_st6_b243_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b243_c0 : nS_st5_b243_c1;
  assign nS_st6_b244_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b244_c0 : nS_st5_b244_c1;
  assign nS_st6_b245_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b245_c0 : nS_st5_b245_c1;
  assign nS_st6_b246_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b246_c0 : nS_st5_b246_c1;
  assign nS_st6_b247_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b247_c0 : nS_st5_b247_c1;
  assign nS_st6_b248_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b248_c0 : nS_st5_b248_c1;
  assign nS_st6_b249_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b249_c0 : nS_st5_b249_c1;
  assign nS_st6_b250_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b250_c0 : nS_st5_b250_c1;
  assign nS_st6_b251_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b251_c0 : nS_st5_b251_c1;
  assign nS_st6_b252_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b252_c0 : nS_st5_b252_c1;
  assign nS_st6_b253_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b253_c0 : nS_st5_b253_c1;
  assign nS_st6_b254_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b254_c0 : nS_st5_b254_c1;
  assign nS_st6_b255_c1 = (nC_st5_b239_c1 == 0) ? nS_st5_b255_c0 : nS_st5_b255_c1;
  assign nC_st6_b31_c0 = (nC_st5_b15_c0 == 0) ? nC_st5_b31_c0 : nC_st5_b31_c1;
  assign nC_st6_b63_c0 = (nC_st5_b47_c0 == 0) ? nC_st5_b63_c0 : nC_st5_b63_c1;
  assign nC_st6_b95_c0 = (nC_st5_b79_c0 == 0) ? nC_st5_b95_c0 : nC_st5_b95_c1;
  assign nC_st6_b127_c0 = (nC_st5_b111_c0 == 0) ? nC_st5_b127_c0 : nC_st5_b127_c1;
  assign nC_st6_b159_c0 = (nC_st5_b143_c0 == 0) ? nC_st5_b159_c0 : nC_st5_b159_c1;
  assign nC_st6_b191_c0 = (nC_st5_b175_c0 == 0) ? nC_st5_b191_c0 : nC_st5_b191_c1;
  assign nC_st6_b223_c0 = (nC_st5_b207_c0 == 0) ? nC_st5_b223_c0 : nC_st5_b223_c1;
  assign nC_st6_b255_c0 = (nC_st5_b239_c0 == 0) ? nC_st5_b255_c0 : nC_st5_b255_c1;
  assign nC_st6_b31_c1 = (nC_st5_b15_c1 == 0) ? nC_st5_b31_c0 : nC_st5_b31_c1;
  assign nC_st6_b63_c1 = (nC_st5_b47_c1 == 0) ? nC_st5_b63_c0 : nC_st5_b63_c1;
  assign nC_st6_b95_c1 = (nC_st5_b79_c1 == 0) ? nC_st5_b95_c0 : nC_st5_b95_c1;
  assign nC_st6_b127_c1 = (nC_st5_b111_c1 == 0) ? nC_st5_b127_c0 : nC_st5_b127_c1;
  assign nC_st6_b159_c1 = (nC_st5_b143_c1 == 0) ? nC_st5_b159_c0 : nC_st5_b159_c1;
  assign nC_st6_b191_c1 = (nC_st5_b175_c1 == 0) ? nC_st5_b191_c0 : nC_st5_b191_c1;
  assign nC_st6_b223_c1 = (nC_st5_b207_c1 == 0) ? nC_st5_b223_c0 : nC_st5_b223_c1;
  assign nC_st6_b255_c1 = (nC_st5_b239_c1 == 0) ? nC_st5_b255_c0 : nC_st5_b255_c1;

  assign nS_st7_b0_c0 = nS_st6_b0_c0;
  assign nS_st7_b1_c0 = nS_st6_b1_c0;
  assign nS_st7_b2_c0 = nS_st6_b2_c0;
  assign nS_st7_b3_c0 = nS_st6_b3_c0;
  assign nS_st7_b4_c0 = nS_st6_b4_c0;
  assign nS_st7_b5_c0 = nS_st6_b5_c0;
  assign nS_st7_b6_c0 = nS_st6_b6_c0;
  assign nS_st7_b7_c0 = nS_st6_b7_c0;
  assign nS_st7_b8_c0 = nS_st6_b8_c0;
  assign nS_st7_b9_c0 = nS_st6_b9_c0;
  assign nS_st7_b10_c0 = nS_st6_b10_c0;
  assign nS_st7_b11_c0 = nS_st6_b11_c0;
  assign nS_st7_b12_c0 = nS_st6_b12_c0;
  assign nS_st7_b13_c0 = nS_st6_b13_c0;
  assign nS_st7_b14_c0 = nS_st6_b14_c0;
  assign nS_st7_b15_c0 = nS_st6_b15_c0;
  assign nS_st7_b16_c0 = nS_st6_b16_c0;
  assign nS_st7_b17_c0 = nS_st6_b17_c0;
  assign nS_st7_b18_c0 = nS_st6_b18_c0;
  assign nS_st7_b19_c0 = nS_st6_b19_c0;
  assign nS_st7_b20_c0 = nS_st6_b20_c0;
  assign nS_st7_b21_c0 = nS_st6_b21_c0;
  assign nS_st7_b22_c0 = nS_st6_b22_c0;
  assign nS_st7_b23_c0 = nS_st6_b23_c0;
  assign nS_st7_b24_c0 = nS_st6_b24_c0;
  assign nS_st7_b25_c0 = nS_st6_b25_c0;
  assign nS_st7_b26_c0 = nS_st6_b26_c0;
  assign nS_st7_b27_c0 = nS_st6_b27_c0;
  assign nS_st7_b28_c0 = nS_st6_b28_c0;
  assign nS_st7_b29_c0 = nS_st6_b29_c0;
  assign nS_st7_b30_c0 = nS_st6_b30_c0;
  assign nS_st7_b31_c0 = nS_st6_b31_c0;
  assign nS_st7_b32_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b32_c0 : nS_st6_b32_c1;
  assign nS_st7_b33_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b33_c0 : nS_st6_b33_c1;
  assign nS_st7_b34_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b34_c0 : nS_st6_b34_c1;
  assign nS_st7_b35_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b35_c0 : nS_st6_b35_c1;
  assign nS_st7_b36_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b36_c0 : nS_st6_b36_c1;
  assign nS_st7_b37_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b37_c0 : nS_st6_b37_c1;
  assign nS_st7_b38_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b38_c0 : nS_st6_b38_c1;
  assign nS_st7_b39_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b39_c0 : nS_st6_b39_c1;
  assign nS_st7_b40_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b40_c0 : nS_st6_b40_c1;
  assign nS_st7_b41_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b41_c0 : nS_st6_b41_c1;
  assign nS_st7_b42_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b42_c0 : nS_st6_b42_c1;
  assign nS_st7_b43_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b43_c0 : nS_st6_b43_c1;
  assign nS_st7_b44_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b44_c0 : nS_st6_b44_c1;
  assign nS_st7_b45_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b45_c0 : nS_st6_b45_c1;
  assign nS_st7_b46_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b46_c0 : nS_st6_b46_c1;
  assign nS_st7_b47_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b47_c0 : nS_st6_b47_c1;
  assign nS_st7_b48_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b48_c0 : nS_st6_b48_c1;
  assign nS_st7_b49_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b49_c0 : nS_st6_b49_c1;
  assign nS_st7_b50_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b50_c0 : nS_st6_b50_c1;
  assign nS_st7_b51_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b51_c0 : nS_st6_b51_c1;
  assign nS_st7_b52_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b52_c0 : nS_st6_b52_c1;
  assign nS_st7_b53_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b53_c0 : nS_st6_b53_c1;
  assign nS_st7_b54_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b54_c0 : nS_st6_b54_c1;
  assign nS_st7_b55_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b55_c0 : nS_st6_b55_c1;
  assign nS_st7_b56_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b56_c0 : nS_st6_b56_c1;
  assign nS_st7_b57_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b57_c0 : nS_st6_b57_c1;
  assign nS_st7_b58_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b58_c0 : nS_st6_b58_c1;
  assign nS_st7_b59_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b59_c0 : nS_st6_b59_c1;
  assign nS_st7_b60_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b60_c0 : nS_st6_b60_c1;
  assign nS_st7_b61_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b61_c0 : nS_st6_b61_c1;
  assign nS_st7_b62_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b62_c0 : nS_st6_b62_c1;
  assign nS_st7_b63_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b63_c0 : nS_st6_b63_c1;
  assign nS_st7_b64_c0 = nS_st6_b64_c0;
  assign nS_st7_b65_c0 = nS_st6_b65_c0;
  assign nS_st7_b66_c0 = nS_st6_b66_c0;
  assign nS_st7_b67_c0 = nS_st6_b67_c0;
  assign nS_st7_b68_c0 = nS_st6_b68_c0;
  assign nS_st7_b69_c0 = nS_st6_b69_c0;
  assign nS_st7_b70_c0 = nS_st6_b70_c0;
  assign nS_st7_b71_c0 = nS_st6_b71_c0;
  assign nS_st7_b72_c0 = nS_st6_b72_c0;
  assign nS_st7_b73_c0 = nS_st6_b73_c0;
  assign nS_st7_b74_c0 = nS_st6_b74_c0;
  assign nS_st7_b75_c0 = nS_st6_b75_c0;
  assign nS_st7_b76_c0 = nS_st6_b76_c0;
  assign nS_st7_b77_c0 = nS_st6_b77_c0;
  assign nS_st7_b78_c0 = nS_st6_b78_c0;
  assign nS_st7_b79_c0 = nS_st6_b79_c0;
  assign nS_st7_b80_c0 = nS_st6_b80_c0;
  assign nS_st7_b81_c0 = nS_st6_b81_c0;
  assign nS_st7_b82_c0 = nS_st6_b82_c0;
  assign nS_st7_b83_c0 = nS_st6_b83_c0;
  assign nS_st7_b84_c0 = nS_st6_b84_c0;
  assign nS_st7_b85_c0 = nS_st6_b85_c0;
  assign nS_st7_b86_c0 = nS_st6_b86_c0;
  assign nS_st7_b87_c0 = nS_st6_b87_c0;
  assign nS_st7_b88_c0 = nS_st6_b88_c0;
  assign nS_st7_b89_c0 = nS_st6_b89_c0;
  assign nS_st7_b90_c0 = nS_st6_b90_c0;
  assign nS_st7_b91_c0 = nS_st6_b91_c0;
  assign nS_st7_b92_c0 = nS_st6_b92_c0;
  assign nS_st7_b93_c0 = nS_st6_b93_c0;
  assign nS_st7_b94_c0 = nS_st6_b94_c0;
  assign nS_st7_b95_c0 = nS_st6_b95_c0;
  assign nS_st7_b96_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b96_c0 : nS_st6_b96_c1;
  assign nS_st7_b97_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b97_c0 : nS_st6_b97_c1;
  assign nS_st7_b98_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b98_c0 : nS_st6_b98_c1;
  assign nS_st7_b99_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b99_c0 : nS_st6_b99_c1;
  assign nS_st7_b100_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b100_c0 : nS_st6_b100_c1;
  assign nS_st7_b101_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b101_c0 : nS_st6_b101_c1;
  assign nS_st7_b102_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b102_c0 : nS_st6_b102_c1;
  assign nS_st7_b103_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b103_c0 : nS_st6_b103_c1;
  assign nS_st7_b104_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b104_c0 : nS_st6_b104_c1;
  assign nS_st7_b105_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b105_c0 : nS_st6_b105_c1;
  assign nS_st7_b106_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b106_c0 : nS_st6_b106_c1;
  assign nS_st7_b107_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b107_c0 : nS_st6_b107_c1;
  assign nS_st7_b108_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b108_c0 : nS_st6_b108_c1;
  assign nS_st7_b109_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b109_c0 : nS_st6_b109_c1;
  assign nS_st7_b110_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b110_c0 : nS_st6_b110_c1;
  assign nS_st7_b111_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b111_c0 : nS_st6_b111_c1;
  assign nS_st7_b112_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b112_c0 : nS_st6_b112_c1;
  assign nS_st7_b113_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b113_c0 : nS_st6_b113_c1;
  assign nS_st7_b114_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b114_c0 : nS_st6_b114_c1;
  assign nS_st7_b115_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b115_c0 : nS_st6_b115_c1;
  assign nS_st7_b116_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b116_c0 : nS_st6_b116_c1;
  assign nS_st7_b117_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b117_c0 : nS_st6_b117_c1;
  assign nS_st7_b118_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b118_c0 : nS_st6_b118_c1;
  assign nS_st7_b119_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b119_c0 : nS_st6_b119_c1;
  assign nS_st7_b120_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b120_c0 : nS_st6_b120_c1;
  assign nS_st7_b121_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b121_c0 : nS_st6_b121_c1;
  assign nS_st7_b122_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b122_c0 : nS_st6_b122_c1;
  assign nS_st7_b123_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b123_c0 : nS_st6_b123_c1;
  assign nS_st7_b124_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b124_c0 : nS_st6_b124_c1;
  assign nS_st7_b125_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b125_c0 : nS_st6_b125_c1;
  assign nS_st7_b126_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b126_c0 : nS_st6_b126_c1;
  assign nS_st7_b127_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b127_c0 : nS_st6_b127_c1;
  assign nS_st7_b128_c0 = nS_st6_b128_c0;
  assign nS_st7_b129_c0 = nS_st6_b129_c0;
  assign nS_st7_b130_c0 = nS_st6_b130_c0;
  assign nS_st7_b131_c0 = nS_st6_b131_c0;
  assign nS_st7_b132_c0 = nS_st6_b132_c0;
  assign nS_st7_b133_c0 = nS_st6_b133_c0;
  assign nS_st7_b134_c0 = nS_st6_b134_c0;
  assign nS_st7_b135_c0 = nS_st6_b135_c0;
  assign nS_st7_b136_c0 = nS_st6_b136_c0;
  assign nS_st7_b137_c0 = nS_st6_b137_c0;
  assign nS_st7_b138_c0 = nS_st6_b138_c0;
  assign nS_st7_b139_c0 = nS_st6_b139_c0;
  assign nS_st7_b140_c0 = nS_st6_b140_c0;
  assign nS_st7_b141_c0 = nS_st6_b141_c0;
  assign nS_st7_b142_c0 = nS_st6_b142_c0;
  assign nS_st7_b143_c0 = nS_st6_b143_c0;
  assign nS_st7_b144_c0 = nS_st6_b144_c0;
  assign nS_st7_b145_c0 = nS_st6_b145_c0;
  assign nS_st7_b146_c0 = nS_st6_b146_c0;
  assign nS_st7_b147_c0 = nS_st6_b147_c0;
  assign nS_st7_b148_c0 = nS_st6_b148_c0;
  assign nS_st7_b149_c0 = nS_st6_b149_c0;
  assign nS_st7_b150_c0 = nS_st6_b150_c0;
  assign nS_st7_b151_c0 = nS_st6_b151_c0;
  assign nS_st7_b152_c0 = nS_st6_b152_c0;
  assign nS_st7_b153_c0 = nS_st6_b153_c0;
  assign nS_st7_b154_c0 = nS_st6_b154_c0;
  assign nS_st7_b155_c0 = nS_st6_b155_c0;
  assign nS_st7_b156_c0 = nS_st6_b156_c0;
  assign nS_st7_b157_c0 = nS_st6_b157_c0;
  assign nS_st7_b158_c0 = nS_st6_b158_c0;
  assign nS_st7_b159_c0 = nS_st6_b159_c0;
  assign nS_st7_b160_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b160_c0 : nS_st6_b160_c1;
  assign nS_st7_b161_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b161_c0 : nS_st6_b161_c1;
  assign nS_st7_b162_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b162_c0 : nS_st6_b162_c1;
  assign nS_st7_b163_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b163_c0 : nS_st6_b163_c1;
  assign nS_st7_b164_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b164_c0 : nS_st6_b164_c1;
  assign nS_st7_b165_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b165_c0 : nS_st6_b165_c1;
  assign nS_st7_b166_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b166_c0 : nS_st6_b166_c1;
  assign nS_st7_b167_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b167_c0 : nS_st6_b167_c1;
  assign nS_st7_b168_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b168_c0 : nS_st6_b168_c1;
  assign nS_st7_b169_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b169_c0 : nS_st6_b169_c1;
  assign nS_st7_b170_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b170_c0 : nS_st6_b170_c1;
  assign nS_st7_b171_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b171_c0 : nS_st6_b171_c1;
  assign nS_st7_b172_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b172_c0 : nS_st6_b172_c1;
  assign nS_st7_b173_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b173_c0 : nS_st6_b173_c1;
  assign nS_st7_b174_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b174_c0 : nS_st6_b174_c1;
  assign nS_st7_b175_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b175_c0 : nS_st6_b175_c1;
  assign nS_st7_b176_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b176_c0 : nS_st6_b176_c1;
  assign nS_st7_b177_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b177_c0 : nS_st6_b177_c1;
  assign nS_st7_b178_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b178_c0 : nS_st6_b178_c1;
  assign nS_st7_b179_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b179_c0 : nS_st6_b179_c1;
  assign nS_st7_b180_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b180_c0 : nS_st6_b180_c1;
  assign nS_st7_b181_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b181_c0 : nS_st6_b181_c1;
  assign nS_st7_b182_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b182_c0 : nS_st6_b182_c1;
  assign nS_st7_b183_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b183_c0 : nS_st6_b183_c1;
  assign nS_st7_b184_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b184_c0 : nS_st6_b184_c1;
  assign nS_st7_b185_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b185_c0 : nS_st6_b185_c1;
  assign nS_st7_b186_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b186_c0 : nS_st6_b186_c1;
  assign nS_st7_b187_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b187_c0 : nS_st6_b187_c1;
  assign nS_st7_b188_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b188_c0 : nS_st6_b188_c1;
  assign nS_st7_b189_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b189_c0 : nS_st6_b189_c1;
  assign nS_st7_b190_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b190_c0 : nS_st6_b190_c1;
  assign nS_st7_b191_c0 = (nC_st6_b159_c0 == 0) ? nS_st6_b191_c0 : nS_st6_b191_c1;
  assign nS_st7_b192_c0 = nS_st6_b192_c0;
  assign nS_st7_b193_c0 = nS_st6_b193_c0;
  assign nS_st7_b194_c0 = nS_st6_b194_c0;
  assign nS_st7_b195_c0 = nS_st6_b195_c0;
  assign nS_st7_b196_c0 = nS_st6_b196_c0;
  assign nS_st7_b197_c0 = nS_st6_b197_c0;
  assign nS_st7_b198_c0 = nS_st6_b198_c0;
  assign nS_st7_b199_c0 = nS_st6_b199_c0;
  assign nS_st7_b200_c0 = nS_st6_b200_c0;
  assign nS_st7_b201_c0 = nS_st6_b201_c0;
  assign nS_st7_b202_c0 = nS_st6_b202_c0;
  assign nS_st7_b203_c0 = nS_st6_b203_c0;
  assign nS_st7_b204_c0 = nS_st6_b204_c0;
  assign nS_st7_b205_c0 = nS_st6_b205_c0;
  assign nS_st7_b206_c0 = nS_st6_b206_c0;
  assign nS_st7_b207_c0 = nS_st6_b207_c0;
  assign nS_st7_b208_c0 = nS_st6_b208_c0;
  assign nS_st7_b209_c0 = nS_st6_b209_c0;
  assign nS_st7_b210_c0 = nS_st6_b210_c0;
  assign nS_st7_b211_c0 = nS_st6_b211_c0;
  assign nS_st7_b212_c0 = nS_st6_b212_c0;
  assign nS_st7_b213_c0 = nS_st6_b213_c0;
  assign nS_st7_b214_c0 = nS_st6_b214_c0;
  assign nS_st7_b215_c0 = nS_st6_b215_c0;
  assign nS_st7_b216_c0 = nS_st6_b216_c0;
  assign nS_st7_b217_c0 = nS_st6_b217_c0;
  assign nS_st7_b218_c0 = nS_st6_b218_c0;
  assign nS_st7_b219_c0 = nS_st6_b219_c0;
  assign nS_st7_b220_c0 = nS_st6_b220_c0;
  assign nS_st7_b221_c0 = nS_st6_b221_c0;
  assign nS_st7_b222_c0 = nS_st6_b222_c0;
  assign nS_st7_b223_c0 = nS_st6_b223_c0;
  assign nS_st7_b224_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b224_c0 : nS_st6_b224_c1;
  assign nS_st7_b225_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b225_c0 : nS_st6_b225_c1;
  assign nS_st7_b226_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b226_c0 : nS_st6_b226_c1;
  assign nS_st7_b227_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b227_c0 : nS_st6_b227_c1;
  assign nS_st7_b228_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b228_c0 : nS_st6_b228_c1;
  assign nS_st7_b229_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b229_c0 : nS_st6_b229_c1;
  assign nS_st7_b230_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b230_c0 : nS_st6_b230_c1;
  assign nS_st7_b231_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b231_c0 : nS_st6_b231_c1;
  assign nS_st7_b232_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b232_c0 : nS_st6_b232_c1;
  assign nS_st7_b233_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b233_c0 : nS_st6_b233_c1;
  assign nS_st7_b234_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b234_c0 : nS_st6_b234_c1;
  assign nS_st7_b235_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b235_c0 : nS_st6_b235_c1;
  assign nS_st7_b236_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b236_c0 : nS_st6_b236_c1;
  assign nS_st7_b237_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b237_c0 : nS_st6_b237_c1;
  assign nS_st7_b238_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b238_c0 : nS_st6_b238_c1;
  assign nS_st7_b239_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b239_c0 : nS_st6_b239_c1;
  assign nS_st7_b240_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b240_c0 : nS_st6_b240_c1;
  assign nS_st7_b241_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b241_c0 : nS_st6_b241_c1;
  assign nS_st7_b242_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b242_c0 : nS_st6_b242_c1;
  assign nS_st7_b243_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b243_c0 : nS_st6_b243_c1;
  assign nS_st7_b244_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b244_c0 : nS_st6_b244_c1;
  assign nS_st7_b245_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b245_c0 : nS_st6_b245_c1;
  assign nS_st7_b246_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b246_c0 : nS_st6_b246_c1;
  assign nS_st7_b247_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b247_c0 : nS_st6_b247_c1;
  assign nS_st7_b248_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b248_c0 : nS_st6_b248_c1;
  assign nS_st7_b249_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b249_c0 : nS_st6_b249_c1;
  assign nS_st7_b250_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b250_c0 : nS_st6_b250_c1;
  assign nS_st7_b251_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b251_c0 : nS_st6_b251_c1;
  assign nS_st7_b252_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b252_c0 : nS_st6_b252_c1;
  assign nS_st7_b253_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b253_c0 : nS_st6_b253_c1;
  assign nS_st7_b254_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b254_c0 : nS_st6_b254_c1;
  assign nS_st7_b255_c0 = (nC_st6_b223_c0 == 0) ? nS_st6_b255_c0 : nS_st6_b255_c1;
  assign nS_st7_b0_c1 = nS_st6_b0_c1;
  assign nS_st7_b1_c1 = nS_st6_b1_c1;
  assign nS_st7_b2_c1 = nS_st6_b2_c1;
  assign nS_st7_b3_c1 = nS_st6_b3_c1;
  assign nS_st7_b4_c1 = nS_st6_b4_c1;
  assign nS_st7_b5_c1 = nS_st6_b5_c1;
  assign nS_st7_b6_c1 = nS_st6_b6_c1;
  assign nS_st7_b7_c1 = nS_st6_b7_c1;
  assign nS_st7_b8_c1 = nS_st6_b8_c1;
  assign nS_st7_b9_c1 = nS_st6_b9_c1;
  assign nS_st7_b10_c1 = nS_st6_b10_c1;
  assign nS_st7_b11_c1 = nS_st6_b11_c1;
  assign nS_st7_b12_c1 = nS_st6_b12_c1;
  assign nS_st7_b13_c1 = nS_st6_b13_c1;
  assign nS_st7_b14_c1 = nS_st6_b14_c1;
  assign nS_st7_b15_c1 = nS_st6_b15_c1;
  assign nS_st7_b16_c1 = nS_st6_b16_c1;
  assign nS_st7_b17_c1 = nS_st6_b17_c1;
  assign nS_st7_b18_c1 = nS_st6_b18_c1;
  assign nS_st7_b19_c1 = nS_st6_b19_c1;
  assign nS_st7_b20_c1 = nS_st6_b20_c1;
  assign nS_st7_b21_c1 = nS_st6_b21_c1;
  assign nS_st7_b22_c1 = nS_st6_b22_c1;
  assign nS_st7_b23_c1 = nS_st6_b23_c1;
  assign nS_st7_b24_c1 = nS_st6_b24_c1;
  assign nS_st7_b25_c1 = nS_st6_b25_c1;
  assign nS_st7_b26_c1 = nS_st6_b26_c1;
  assign nS_st7_b27_c1 = nS_st6_b27_c1;
  assign nS_st7_b28_c1 = nS_st6_b28_c1;
  assign nS_st7_b29_c1 = nS_st6_b29_c1;
  assign nS_st7_b30_c1 = nS_st6_b30_c1;
  assign nS_st7_b31_c1 = nS_st6_b31_c1;
  assign nS_st7_b32_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b32_c0 : nS_st6_b32_c1;
  assign nS_st7_b33_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b33_c0 : nS_st6_b33_c1;
  assign nS_st7_b34_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b34_c0 : nS_st6_b34_c1;
  assign nS_st7_b35_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b35_c0 : nS_st6_b35_c1;
  assign nS_st7_b36_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b36_c0 : nS_st6_b36_c1;
  assign nS_st7_b37_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b37_c0 : nS_st6_b37_c1;
  assign nS_st7_b38_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b38_c0 : nS_st6_b38_c1;
  assign nS_st7_b39_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b39_c0 : nS_st6_b39_c1;
  assign nS_st7_b40_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b40_c0 : nS_st6_b40_c1;
  assign nS_st7_b41_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b41_c0 : nS_st6_b41_c1;
  assign nS_st7_b42_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b42_c0 : nS_st6_b42_c1;
  assign nS_st7_b43_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b43_c0 : nS_st6_b43_c1;
  assign nS_st7_b44_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b44_c0 : nS_st6_b44_c1;
  assign nS_st7_b45_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b45_c0 : nS_st6_b45_c1;
  assign nS_st7_b46_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b46_c0 : nS_st6_b46_c1;
  assign nS_st7_b47_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b47_c0 : nS_st6_b47_c1;
  assign nS_st7_b48_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b48_c0 : nS_st6_b48_c1;
  assign nS_st7_b49_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b49_c0 : nS_st6_b49_c1;
  assign nS_st7_b50_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b50_c0 : nS_st6_b50_c1;
  assign nS_st7_b51_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b51_c0 : nS_st6_b51_c1;
  assign nS_st7_b52_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b52_c0 : nS_st6_b52_c1;
  assign nS_st7_b53_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b53_c0 : nS_st6_b53_c1;
  assign nS_st7_b54_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b54_c0 : nS_st6_b54_c1;
  assign nS_st7_b55_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b55_c0 : nS_st6_b55_c1;
  assign nS_st7_b56_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b56_c0 : nS_st6_b56_c1;
  assign nS_st7_b57_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b57_c0 : nS_st6_b57_c1;
  assign nS_st7_b58_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b58_c0 : nS_st6_b58_c1;
  assign nS_st7_b59_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b59_c0 : nS_st6_b59_c1;
  assign nS_st7_b60_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b60_c0 : nS_st6_b60_c1;
  assign nS_st7_b61_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b61_c0 : nS_st6_b61_c1;
  assign nS_st7_b62_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b62_c0 : nS_st6_b62_c1;
  assign nS_st7_b63_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b63_c0 : nS_st6_b63_c1;
  assign nS_st7_b64_c1 = nS_st6_b64_c1;
  assign nS_st7_b65_c1 = nS_st6_b65_c1;
  assign nS_st7_b66_c1 = nS_st6_b66_c1;
  assign nS_st7_b67_c1 = nS_st6_b67_c1;
  assign nS_st7_b68_c1 = nS_st6_b68_c1;
  assign nS_st7_b69_c1 = nS_st6_b69_c1;
  assign nS_st7_b70_c1 = nS_st6_b70_c1;
  assign nS_st7_b71_c1 = nS_st6_b71_c1;
  assign nS_st7_b72_c1 = nS_st6_b72_c1;
  assign nS_st7_b73_c1 = nS_st6_b73_c1;
  assign nS_st7_b74_c1 = nS_st6_b74_c1;
  assign nS_st7_b75_c1 = nS_st6_b75_c1;
  assign nS_st7_b76_c1 = nS_st6_b76_c1;
  assign nS_st7_b77_c1 = nS_st6_b77_c1;
  assign nS_st7_b78_c1 = nS_st6_b78_c1;
  assign nS_st7_b79_c1 = nS_st6_b79_c1;
  assign nS_st7_b80_c1 = nS_st6_b80_c1;
  assign nS_st7_b81_c1 = nS_st6_b81_c1;
  assign nS_st7_b82_c1 = nS_st6_b82_c1;
  assign nS_st7_b83_c1 = nS_st6_b83_c1;
  assign nS_st7_b84_c1 = nS_st6_b84_c1;
  assign nS_st7_b85_c1 = nS_st6_b85_c1;
  assign nS_st7_b86_c1 = nS_st6_b86_c1;
  assign nS_st7_b87_c1 = nS_st6_b87_c1;
  assign nS_st7_b88_c1 = nS_st6_b88_c1;
  assign nS_st7_b89_c1 = nS_st6_b89_c1;
  assign nS_st7_b90_c1 = nS_st6_b90_c1;
  assign nS_st7_b91_c1 = nS_st6_b91_c1;
  assign nS_st7_b92_c1 = nS_st6_b92_c1;
  assign nS_st7_b93_c1 = nS_st6_b93_c1;
  assign nS_st7_b94_c1 = nS_st6_b94_c1;
  assign nS_st7_b95_c1 = nS_st6_b95_c1;
  assign nS_st7_b96_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b96_c0 : nS_st6_b96_c1;
  assign nS_st7_b97_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b97_c0 : nS_st6_b97_c1;
  assign nS_st7_b98_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b98_c0 : nS_st6_b98_c1;
  assign nS_st7_b99_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b99_c0 : nS_st6_b99_c1;
  assign nS_st7_b100_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b100_c0 : nS_st6_b100_c1;
  assign nS_st7_b101_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b101_c0 : nS_st6_b101_c1;
  assign nS_st7_b102_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b102_c0 : nS_st6_b102_c1;
  assign nS_st7_b103_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b103_c0 : nS_st6_b103_c1;
  assign nS_st7_b104_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b104_c0 : nS_st6_b104_c1;
  assign nS_st7_b105_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b105_c0 : nS_st6_b105_c1;
  assign nS_st7_b106_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b106_c0 : nS_st6_b106_c1;
  assign nS_st7_b107_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b107_c0 : nS_st6_b107_c1;
  assign nS_st7_b108_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b108_c0 : nS_st6_b108_c1;
  assign nS_st7_b109_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b109_c0 : nS_st6_b109_c1;
  assign nS_st7_b110_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b110_c0 : nS_st6_b110_c1;
  assign nS_st7_b111_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b111_c0 : nS_st6_b111_c1;
  assign nS_st7_b112_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b112_c0 : nS_st6_b112_c1;
  assign nS_st7_b113_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b113_c0 : nS_st6_b113_c1;
  assign nS_st7_b114_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b114_c0 : nS_st6_b114_c1;
  assign nS_st7_b115_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b115_c0 : nS_st6_b115_c1;
  assign nS_st7_b116_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b116_c0 : nS_st6_b116_c1;
  assign nS_st7_b117_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b117_c0 : nS_st6_b117_c1;
  assign nS_st7_b118_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b118_c0 : nS_st6_b118_c1;
  assign nS_st7_b119_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b119_c0 : nS_st6_b119_c1;
  assign nS_st7_b120_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b120_c0 : nS_st6_b120_c1;
  assign nS_st7_b121_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b121_c0 : nS_st6_b121_c1;
  assign nS_st7_b122_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b122_c0 : nS_st6_b122_c1;
  assign nS_st7_b123_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b123_c0 : nS_st6_b123_c1;
  assign nS_st7_b124_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b124_c0 : nS_st6_b124_c1;
  assign nS_st7_b125_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b125_c0 : nS_st6_b125_c1;
  assign nS_st7_b126_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b126_c0 : nS_st6_b126_c1;
  assign nS_st7_b127_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b127_c0 : nS_st6_b127_c1;
  assign nS_st7_b128_c1 = nS_st6_b128_c1;
  assign nS_st7_b129_c1 = nS_st6_b129_c1;
  assign nS_st7_b130_c1 = nS_st6_b130_c1;
  assign nS_st7_b131_c1 = nS_st6_b131_c1;
  assign nS_st7_b132_c1 = nS_st6_b132_c1;
  assign nS_st7_b133_c1 = nS_st6_b133_c1;
  assign nS_st7_b134_c1 = nS_st6_b134_c1;
  assign nS_st7_b135_c1 = nS_st6_b135_c1;
  assign nS_st7_b136_c1 = nS_st6_b136_c1;
  assign nS_st7_b137_c1 = nS_st6_b137_c1;
  assign nS_st7_b138_c1 = nS_st6_b138_c1;
  assign nS_st7_b139_c1 = nS_st6_b139_c1;
  assign nS_st7_b140_c1 = nS_st6_b140_c1;
  assign nS_st7_b141_c1 = nS_st6_b141_c1;
  assign nS_st7_b142_c1 = nS_st6_b142_c1;
  assign nS_st7_b143_c1 = nS_st6_b143_c1;
  assign nS_st7_b144_c1 = nS_st6_b144_c1;
  assign nS_st7_b145_c1 = nS_st6_b145_c1;
  assign nS_st7_b146_c1 = nS_st6_b146_c1;
  assign nS_st7_b147_c1 = nS_st6_b147_c1;
  assign nS_st7_b148_c1 = nS_st6_b148_c1;
  assign nS_st7_b149_c1 = nS_st6_b149_c1;
  assign nS_st7_b150_c1 = nS_st6_b150_c1;
  assign nS_st7_b151_c1 = nS_st6_b151_c1;
  assign nS_st7_b152_c1 = nS_st6_b152_c1;
  assign nS_st7_b153_c1 = nS_st6_b153_c1;
  assign nS_st7_b154_c1 = nS_st6_b154_c1;
  assign nS_st7_b155_c1 = nS_st6_b155_c1;
  assign nS_st7_b156_c1 = nS_st6_b156_c1;
  assign nS_st7_b157_c1 = nS_st6_b157_c1;
  assign nS_st7_b158_c1 = nS_st6_b158_c1;
  assign nS_st7_b159_c1 = nS_st6_b159_c1;
  assign nS_st7_b160_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b160_c0 : nS_st6_b160_c1;
  assign nS_st7_b161_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b161_c0 : nS_st6_b161_c1;
  assign nS_st7_b162_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b162_c0 : nS_st6_b162_c1;
  assign nS_st7_b163_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b163_c0 : nS_st6_b163_c1;
  assign nS_st7_b164_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b164_c0 : nS_st6_b164_c1;
  assign nS_st7_b165_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b165_c0 : nS_st6_b165_c1;
  assign nS_st7_b166_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b166_c0 : nS_st6_b166_c1;
  assign nS_st7_b167_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b167_c0 : nS_st6_b167_c1;
  assign nS_st7_b168_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b168_c0 : nS_st6_b168_c1;
  assign nS_st7_b169_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b169_c0 : nS_st6_b169_c1;
  assign nS_st7_b170_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b170_c0 : nS_st6_b170_c1;
  assign nS_st7_b171_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b171_c0 : nS_st6_b171_c1;
  assign nS_st7_b172_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b172_c0 : nS_st6_b172_c1;
  assign nS_st7_b173_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b173_c0 : nS_st6_b173_c1;
  assign nS_st7_b174_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b174_c0 : nS_st6_b174_c1;
  assign nS_st7_b175_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b175_c0 : nS_st6_b175_c1;
  assign nS_st7_b176_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b176_c0 : nS_st6_b176_c1;
  assign nS_st7_b177_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b177_c0 : nS_st6_b177_c1;
  assign nS_st7_b178_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b178_c0 : nS_st6_b178_c1;
  assign nS_st7_b179_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b179_c0 : nS_st6_b179_c1;
  assign nS_st7_b180_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b180_c0 : nS_st6_b180_c1;
  assign nS_st7_b181_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b181_c0 : nS_st6_b181_c1;
  assign nS_st7_b182_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b182_c0 : nS_st6_b182_c1;
  assign nS_st7_b183_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b183_c0 : nS_st6_b183_c1;
  assign nS_st7_b184_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b184_c0 : nS_st6_b184_c1;
  assign nS_st7_b185_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b185_c0 : nS_st6_b185_c1;
  assign nS_st7_b186_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b186_c0 : nS_st6_b186_c1;
  assign nS_st7_b187_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b187_c0 : nS_st6_b187_c1;
  assign nS_st7_b188_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b188_c0 : nS_st6_b188_c1;
  assign nS_st7_b189_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b189_c0 : nS_st6_b189_c1;
  assign nS_st7_b190_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b190_c0 : nS_st6_b190_c1;
  assign nS_st7_b191_c1 = (nC_st6_b159_c1 == 0) ? nS_st6_b191_c0 : nS_st6_b191_c1;
  assign nS_st7_b192_c1 = nS_st6_b192_c1;
  assign nS_st7_b193_c1 = nS_st6_b193_c1;
  assign nS_st7_b194_c1 = nS_st6_b194_c1;
  assign nS_st7_b195_c1 = nS_st6_b195_c1;
  assign nS_st7_b196_c1 = nS_st6_b196_c1;
  assign nS_st7_b197_c1 = nS_st6_b197_c1;
  assign nS_st7_b198_c1 = nS_st6_b198_c1;
  assign nS_st7_b199_c1 = nS_st6_b199_c1;
  assign nS_st7_b200_c1 = nS_st6_b200_c1;
  assign nS_st7_b201_c1 = nS_st6_b201_c1;
  assign nS_st7_b202_c1 = nS_st6_b202_c1;
  assign nS_st7_b203_c1 = nS_st6_b203_c1;
  assign nS_st7_b204_c1 = nS_st6_b204_c1;
  assign nS_st7_b205_c1 = nS_st6_b205_c1;
  assign nS_st7_b206_c1 = nS_st6_b206_c1;
  assign nS_st7_b207_c1 = nS_st6_b207_c1;
  assign nS_st7_b208_c1 = nS_st6_b208_c1;
  assign nS_st7_b209_c1 = nS_st6_b209_c1;
  assign nS_st7_b210_c1 = nS_st6_b210_c1;
  assign nS_st7_b211_c1 = nS_st6_b211_c1;
  assign nS_st7_b212_c1 = nS_st6_b212_c1;
  assign nS_st7_b213_c1 = nS_st6_b213_c1;
  assign nS_st7_b214_c1 = nS_st6_b214_c1;
  assign nS_st7_b215_c1 = nS_st6_b215_c1;
  assign nS_st7_b216_c1 = nS_st6_b216_c1;
  assign nS_st7_b217_c1 = nS_st6_b217_c1;
  assign nS_st7_b218_c1 = nS_st6_b218_c1;
  assign nS_st7_b219_c1 = nS_st6_b219_c1;
  assign nS_st7_b220_c1 = nS_st6_b220_c1;
  assign nS_st7_b221_c1 = nS_st6_b221_c1;
  assign nS_st7_b222_c1 = nS_st6_b222_c1;
  assign nS_st7_b223_c1 = nS_st6_b223_c1;
  assign nS_st7_b224_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b224_c0 : nS_st6_b224_c1;
  assign nS_st7_b225_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b225_c0 : nS_st6_b225_c1;
  assign nS_st7_b226_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b226_c0 : nS_st6_b226_c1;
  assign nS_st7_b227_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b227_c0 : nS_st6_b227_c1;
  assign nS_st7_b228_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b228_c0 : nS_st6_b228_c1;
  assign nS_st7_b229_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b229_c0 : nS_st6_b229_c1;
  assign nS_st7_b230_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b230_c0 : nS_st6_b230_c1;
  assign nS_st7_b231_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b231_c0 : nS_st6_b231_c1;
  assign nS_st7_b232_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b232_c0 : nS_st6_b232_c1;
  assign nS_st7_b233_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b233_c0 : nS_st6_b233_c1;
  assign nS_st7_b234_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b234_c0 : nS_st6_b234_c1;
  assign nS_st7_b235_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b235_c0 : nS_st6_b235_c1;
  assign nS_st7_b236_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b236_c0 : nS_st6_b236_c1;
  assign nS_st7_b237_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b237_c0 : nS_st6_b237_c1;
  assign nS_st7_b238_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b238_c0 : nS_st6_b238_c1;
  assign nS_st7_b239_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b239_c0 : nS_st6_b239_c1;
  assign nS_st7_b240_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b240_c0 : nS_st6_b240_c1;
  assign nS_st7_b241_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b241_c0 : nS_st6_b241_c1;
  assign nS_st7_b242_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b242_c0 : nS_st6_b242_c1;
  assign nS_st7_b243_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b243_c0 : nS_st6_b243_c1;
  assign nS_st7_b244_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b244_c0 : nS_st6_b244_c1;
  assign nS_st7_b245_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b245_c0 : nS_st6_b245_c1;
  assign nS_st7_b246_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b246_c0 : nS_st6_b246_c1;
  assign nS_st7_b247_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b247_c0 : nS_st6_b247_c1;
  assign nS_st7_b248_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b248_c0 : nS_st6_b248_c1;
  assign nS_st7_b249_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b249_c0 : nS_st6_b249_c1;
  assign nS_st7_b250_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b250_c0 : nS_st6_b250_c1;
  assign nS_st7_b251_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b251_c0 : nS_st6_b251_c1;
  assign nS_st7_b252_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b252_c0 : nS_st6_b252_c1;
  assign nS_st7_b253_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b253_c0 : nS_st6_b253_c1;
  assign nS_st7_b254_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b254_c0 : nS_st6_b254_c1;
  assign nS_st7_b255_c1 = (nC_st6_b223_c1 == 0) ? nS_st6_b255_c0 : nS_st6_b255_c1;
  assign nC_st7_b63_c0 = (nC_st6_b31_c0 == 0) ? nC_st6_b63_c0 : nC_st6_b63_c1;
  assign nC_st7_b127_c0 = (nC_st6_b95_c0 == 0) ? nC_st6_b127_c0 : nC_st6_b127_c1;
  assign nC_st7_b191_c0 = (nC_st6_b159_c0 == 0) ? nC_st6_b191_c0 : nC_st6_b191_c1;
  assign nC_st7_b255_c0 = (nC_st6_b223_c0 == 0) ? nC_st6_b255_c0 : nC_st6_b255_c1;
  assign nC_st7_b63_c1 = (nC_st6_b31_c1 == 0) ? nC_st6_b63_c0 : nC_st6_b63_c1;
  assign nC_st7_b127_c1 = (nC_st6_b95_c1 == 0) ? nC_st6_b127_c0 : nC_st6_b127_c1;
  assign nC_st7_b191_c1 = (nC_st6_b159_c1 == 0) ? nC_st6_b191_c0 : nC_st6_b191_c1;
  assign nC_st7_b255_c1 = (nC_st6_b223_c1 == 0) ? nC_st6_b255_c0 : nC_st6_b255_c1;

  assign nS_st8_b0_c0 = nS_st7_b0_c0;
  assign nS_st8_b1_c0 = nS_st7_b1_c0;
  assign nS_st8_b2_c0 = nS_st7_b2_c0;
  assign nS_st8_b3_c0 = nS_st7_b3_c0;
  assign nS_st8_b4_c0 = nS_st7_b4_c0;
  assign nS_st8_b5_c0 = nS_st7_b5_c0;
  assign nS_st8_b6_c0 = nS_st7_b6_c0;
  assign nS_st8_b7_c0 = nS_st7_b7_c0;
  assign nS_st8_b8_c0 = nS_st7_b8_c0;
  assign nS_st8_b9_c0 = nS_st7_b9_c0;
  assign nS_st8_b10_c0 = nS_st7_b10_c0;
  assign nS_st8_b11_c0 = nS_st7_b11_c0;
  assign nS_st8_b12_c0 = nS_st7_b12_c0;
  assign nS_st8_b13_c0 = nS_st7_b13_c0;
  assign nS_st8_b14_c0 = nS_st7_b14_c0;
  assign nS_st8_b15_c0 = nS_st7_b15_c0;
  assign nS_st8_b16_c0 = nS_st7_b16_c0;
  assign nS_st8_b17_c0 = nS_st7_b17_c0;
  assign nS_st8_b18_c0 = nS_st7_b18_c0;
  assign nS_st8_b19_c0 = nS_st7_b19_c0;
  assign nS_st8_b20_c0 = nS_st7_b20_c0;
  assign nS_st8_b21_c0 = nS_st7_b21_c0;
  assign nS_st8_b22_c0 = nS_st7_b22_c0;
  assign nS_st8_b23_c0 = nS_st7_b23_c0;
  assign nS_st8_b24_c0 = nS_st7_b24_c0;
  assign nS_st8_b25_c0 = nS_st7_b25_c0;
  assign nS_st8_b26_c0 = nS_st7_b26_c0;
  assign nS_st8_b27_c0 = nS_st7_b27_c0;
  assign nS_st8_b28_c0 = nS_st7_b28_c0;
  assign nS_st8_b29_c0 = nS_st7_b29_c0;
  assign nS_st8_b30_c0 = nS_st7_b30_c0;
  assign nS_st8_b31_c0 = nS_st7_b31_c0;
  assign nS_st8_b32_c0 = nS_st7_b32_c0;
  assign nS_st8_b33_c0 = nS_st7_b33_c0;
  assign nS_st8_b34_c0 = nS_st7_b34_c0;
  assign nS_st8_b35_c0 = nS_st7_b35_c0;
  assign nS_st8_b36_c0 = nS_st7_b36_c0;
  assign nS_st8_b37_c0 = nS_st7_b37_c0;
  assign nS_st8_b38_c0 = nS_st7_b38_c0;
  assign nS_st8_b39_c0 = nS_st7_b39_c0;
  assign nS_st8_b40_c0 = nS_st7_b40_c0;
  assign nS_st8_b41_c0 = nS_st7_b41_c0;
  assign nS_st8_b42_c0 = nS_st7_b42_c0;
  assign nS_st8_b43_c0 = nS_st7_b43_c0;
  assign nS_st8_b44_c0 = nS_st7_b44_c0;
  assign nS_st8_b45_c0 = nS_st7_b45_c0;
  assign nS_st8_b46_c0 = nS_st7_b46_c0;
  assign nS_st8_b47_c0 = nS_st7_b47_c0;
  assign nS_st8_b48_c0 = nS_st7_b48_c0;
  assign nS_st8_b49_c0 = nS_st7_b49_c0;
  assign nS_st8_b50_c0 = nS_st7_b50_c0;
  assign nS_st8_b51_c0 = nS_st7_b51_c0;
  assign nS_st8_b52_c0 = nS_st7_b52_c0;
  assign nS_st8_b53_c0 = nS_st7_b53_c0;
  assign nS_st8_b54_c0 = nS_st7_b54_c0;
  assign nS_st8_b55_c0 = nS_st7_b55_c0;
  assign nS_st8_b56_c0 = nS_st7_b56_c0;
  assign nS_st8_b57_c0 = nS_st7_b57_c0;
  assign nS_st8_b58_c0 = nS_st7_b58_c0;
  assign nS_st8_b59_c0 = nS_st7_b59_c0;
  assign nS_st8_b60_c0 = nS_st7_b60_c0;
  assign nS_st8_b61_c0 = nS_st7_b61_c0;
  assign nS_st8_b62_c0 = nS_st7_b62_c0;
  assign nS_st8_b63_c0 = nS_st7_b63_c0;
  assign nS_st8_b64_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b64_c0 : nS_st7_b64_c1;
  assign nS_st8_b65_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b65_c0 : nS_st7_b65_c1;
  assign nS_st8_b66_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b66_c0 : nS_st7_b66_c1;
  assign nS_st8_b67_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b67_c0 : nS_st7_b67_c1;
  assign nS_st8_b68_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b68_c0 : nS_st7_b68_c1;
  assign nS_st8_b69_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b69_c0 : nS_st7_b69_c1;
  assign nS_st8_b70_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b70_c0 : nS_st7_b70_c1;
  assign nS_st8_b71_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b71_c0 : nS_st7_b71_c1;
  assign nS_st8_b72_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b72_c0 : nS_st7_b72_c1;
  assign nS_st8_b73_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b73_c0 : nS_st7_b73_c1;
  assign nS_st8_b74_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b74_c0 : nS_st7_b74_c1;
  assign nS_st8_b75_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b75_c0 : nS_st7_b75_c1;
  assign nS_st8_b76_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b76_c0 : nS_st7_b76_c1;
  assign nS_st8_b77_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b77_c0 : nS_st7_b77_c1;
  assign nS_st8_b78_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b78_c0 : nS_st7_b78_c1;
  assign nS_st8_b79_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b79_c0 : nS_st7_b79_c1;
  assign nS_st8_b80_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b80_c0 : nS_st7_b80_c1;
  assign nS_st8_b81_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b81_c0 : nS_st7_b81_c1;
  assign nS_st8_b82_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b82_c0 : nS_st7_b82_c1;
  assign nS_st8_b83_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b83_c0 : nS_st7_b83_c1;
  assign nS_st8_b84_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b84_c0 : nS_st7_b84_c1;
  assign nS_st8_b85_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b85_c0 : nS_st7_b85_c1;
  assign nS_st8_b86_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b86_c0 : nS_st7_b86_c1;
  assign nS_st8_b87_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b87_c0 : nS_st7_b87_c1;
  assign nS_st8_b88_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b88_c0 : nS_st7_b88_c1;
  assign nS_st8_b89_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b89_c0 : nS_st7_b89_c1;
  assign nS_st8_b90_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b90_c0 : nS_st7_b90_c1;
  assign nS_st8_b91_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b91_c0 : nS_st7_b91_c1;
  assign nS_st8_b92_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b92_c0 : nS_st7_b92_c1;
  assign nS_st8_b93_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b93_c0 : nS_st7_b93_c1;
  assign nS_st8_b94_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b94_c0 : nS_st7_b94_c1;
  assign nS_st8_b95_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b95_c0 : nS_st7_b95_c1;
  assign nS_st8_b96_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b96_c0 : nS_st7_b96_c1;
  assign nS_st8_b97_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b97_c0 : nS_st7_b97_c1;
  assign nS_st8_b98_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b98_c0 : nS_st7_b98_c1;
  assign nS_st8_b99_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b99_c0 : nS_st7_b99_c1;
  assign nS_st8_b100_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b100_c0 : nS_st7_b100_c1;
  assign nS_st8_b101_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b101_c0 : nS_st7_b101_c1;
  assign nS_st8_b102_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b102_c0 : nS_st7_b102_c1;
  assign nS_st8_b103_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b103_c0 : nS_st7_b103_c1;
  assign nS_st8_b104_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b104_c0 : nS_st7_b104_c1;
  assign nS_st8_b105_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b105_c0 : nS_st7_b105_c1;
  assign nS_st8_b106_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b106_c0 : nS_st7_b106_c1;
  assign nS_st8_b107_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b107_c0 : nS_st7_b107_c1;
  assign nS_st8_b108_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b108_c0 : nS_st7_b108_c1;
  assign nS_st8_b109_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b109_c0 : nS_st7_b109_c1;
  assign nS_st8_b110_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b110_c0 : nS_st7_b110_c1;
  assign nS_st8_b111_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b111_c0 : nS_st7_b111_c1;
  assign nS_st8_b112_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b112_c0 : nS_st7_b112_c1;
  assign nS_st8_b113_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b113_c0 : nS_st7_b113_c1;
  assign nS_st8_b114_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b114_c0 : nS_st7_b114_c1;
  assign nS_st8_b115_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b115_c0 : nS_st7_b115_c1;
  assign nS_st8_b116_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b116_c0 : nS_st7_b116_c1;
  assign nS_st8_b117_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b117_c0 : nS_st7_b117_c1;
  assign nS_st8_b118_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b118_c0 : nS_st7_b118_c1;
  assign nS_st8_b119_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b119_c0 : nS_st7_b119_c1;
  assign nS_st8_b120_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b120_c0 : nS_st7_b120_c1;
  assign nS_st8_b121_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b121_c0 : nS_st7_b121_c1;
  assign nS_st8_b122_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b122_c0 : nS_st7_b122_c1;
  assign nS_st8_b123_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b123_c0 : nS_st7_b123_c1;
  assign nS_st8_b124_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b124_c0 : nS_st7_b124_c1;
  assign nS_st8_b125_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b125_c0 : nS_st7_b125_c1;
  assign nS_st8_b126_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b126_c0 : nS_st7_b126_c1;
  assign nS_st8_b127_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b127_c0 : nS_st7_b127_c1;
  assign nS_st8_b128_c0 = nS_st7_b128_c0;
  assign nS_st8_b129_c0 = nS_st7_b129_c0;
  assign nS_st8_b130_c0 = nS_st7_b130_c0;
  assign nS_st8_b131_c0 = nS_st7_b131_c0;
  assign nS_st8_b132_c0 = nS_st7_b132_c0;
  assign nS_st8_b133_c0 = nS_st7_b133_c0;
  assign nS_st8_b134_c0 = nS_st7_b134_c0;
  assign nS_st8_b135_c0 = nS_st7_b135_c0;
  assign nS_st8_b136_c0 = nS_st7_b136_c0;
  assign nS_st8_b137_c0 = nS_st7_b137_c0;
  assign nS_st8_b138_c0 = nS_st7_b138_c0;
  assign nS_st8_b139_c0 = nS_st7_b139_c0;
  assign nS_st8_b140_c0 = nS_st7_b140_c0;
  assign nS_st8_b141_c0 = nS_st7_b141_c0;
  assign nS_st8_b142_c0 = nS_st7_b142_c0;
  assign nS_st8_b143_c0 = nS_st7_b143_c0;
  assign nS_st8_b144_c0 = nS_st7_b144_c0;
  assign nS_st8_b145_c0 = nS_st7_b145_c0;
  assign nS_st8_b146_c0 = nS_st7_b146_c0;
  assign nS_st8_b147_c0 = nS_st7_b147_c0;
  assign nS_st8_b148_c0 = nS_st7_b148_c0;
  assign nS_st8_b149_c0 = nS_st7_b149_c0;
  assign nS_st8_b150_c0 = nS_st7_b150_c0;
  assign nS_st8_b151_c0 = nS_st7_b151_c0;
  assign nS_st8_b152_c0 = nS_st7_b152_c0;
  assign nS_st8_b153_c0 = nS_st7_b153_c0;
  assign nS_st8_b154_c0 = nS_st7_b154_c0;
  assign nS_st8_b155_c0 = nS_st7_b155_c0;
  assign nS_st8_b156_c0 = nS_st7_b156_c0;
  assign nS_st8_b157_c0 = nS_st7_b157_c0;
  assign nS_st8_b158_c0 = nS_st7_b158_c0;
  assign nS_st8_b159_c0 = nS_st7_b159_c0;
  assign nS_st8_b160_c0 = nS_st7_b160_c0;
  assign nS_st8_b161_c0 = nS_st7_b161_c0;
  assign nS_st8_b162_c0 = nS_st7_b162_c0;
  assign nS_st8_b163_c0 = nS_st7_b163_c0;
  assign nS_st8_b164_c0 = nS_st7_b164_c0;
  assign nS_st8_b165_c0 = nS_st7_b165_c0;
  assign nS_st8_b166_c0 = nS_st7_b166_c0;
  assign nS_st8_b167_c0 = nS_st7_b167_c0;
  assign nS_st8_b168_c0 = nS_st7_b168_c0;
  assign nS_st8_b169_c0 = nS_st7_b169_c0;
  assign nS_st8_b170_c0 = nS_st7_b170_c0;
  assign nS_st8_b171_c0 = nS_st7_b171_c0;
  assign nS_st8_b172_c0 = nS_st7_b172_c0;
  assign nS_st8_b173_c0 = nS_st7_b173_c0;
  assign nS_st8_b174_c0 = nS_st7_b174_c0;
  assign nS_st8_b175_c0 = nS_st7_b175_c0;
  assign nS_st8_b176_c0 = nS_st7_b176_c0;
  assign nS_st8_b177_c0 = nS_st7_b177_c0;
  assign nS_st8_b178_c0 = nS_st7_b178_c0;
  assign nS_st8_b179_c0 = nS_st7_b179_c0;
  assign nS_st8_b180_c0 = nS_st7_b180_c0;
  assign nS_st8_b181_c0 = nS_st7_b181_c0;
  assign nS_st8_b182_c0 = nS_st7_b182_c0;
  assign nS_st8_b183_c0 = nS_st7_b183_c0;
  assign nS_st8_b184_c0 = nS_st7_b184_c0;
  assign nS_st8_b185_c0 = nS_st7_b185_c0;
  assign nS_st8_b186_c0 = nS_st7_b186_c0;
  assign nS_st8_b187_c0 = nS_st7_b187_c0;
  assign nS_st8_b188_c0 = nS_st7_b188_c0;
  assign nS_st8_b189_c0 = nS_st7_b189_c0;
  assign nS_st8_b190_c0 = nS_st7_b190_c0;
  assign nS_st8_b191_c0 = nS_st7_b191_c0;
  assign nS_st8_b192_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b192_c0 : nS_st7_b192_c1;
  assign nS_st8_b193_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b193_c0 : nS_st7_b193_c1;
  assign nS_st8_b194_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b194_c0 : nS_st7_b194_c1;
  assign nS_st8_b195_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b195_c0 : nS_st7_b195_c1;
  assign nS_st8_b196_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b196_c0 : nS_st7_b196_c1;
  assign nS_st8_b197_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b197_c0 : nS_st7_b197_c1;
  assign nS_st8_b198_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b198_c0 : nS_st7_b198_c1;
  assign nS_st8_b199_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b199_c0 : nS_st7_b199_c1;
  assign nS_st8_b200_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b200_c0 : nS_st7_b200_c1;
  assign nS_st8_b201_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b201_c0 : nS_st7_b201_c1;
  assign nS_st8_b202_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b202_c0 : nS_st7_b202_c1;
  assign nS_st8_b203_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b203_c0 : nS_st7_b203_c1;
  assign nS_st8_b204_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b204_c0 : nS_st7_b204_c1;
  assign nS_st8_b205_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b205_c0 : nS_st7_b205_c1;
  assign nS_st8_b206_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b206_c0 : nS_st7_b206_c1;
  assign nS_st8_b207_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b207_c0 : nS_st7_b207_c1;
  assign nS_st8_b208_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b208_c0 : nS_st7_b208_c1;
  assign nS_st8_b209_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b209_c0 : nS_st7_b209_c1;
  assign nS_st8_b210_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b210_c0 : nS_st7_b210_c1;
  assign nS_st8_b211_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b211_c0 : nS_st7_b211_c1;
  assign nS_st8_b212_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b212_c0 : nS_st7_b212_c1;
  assign nS_st8_b213_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b213_c0 : nS_st7_b213_c1;
  assign nS_st8_b214_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b214_c0 : nS_st7_b214_c1;
  assign nS_st8_b215_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b215_c0 : nS_st7_b215_c1;
  assign nS_st8_b216_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b216_c0 : nS_st7_b216_c1;
  assign nS_st8_b217_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b217_c0 : nS_st7_b217_c1;
  assign nS_st8_b218_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b218_c0 : nS_st7_b218_c1;
  assign nS_st8_b219_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b219_c0 : nS_st7_b219_c1;
  assign nS_st8_b220_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b220_c0 : nS_st7_b220_c1;
  assign nS_st8_b221_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b221_c0 : nS_st7_b221_c1;
  assign nS_st8_b222_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b222_c0 : nS_st7_b222_c1;
  assign nS_st8_b223_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b223_c0 : nS_st7_b223_c1;
  assign nS_st8_b224_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b224_c0 : nS_st7_b224_c1;
  assign nS_st8_b225_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b225_c0 : nS_st7_b225_c1;
  assign nS_st8_b226_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b226_c0 : nS_st7_b226_c1;
  assign nS_st8_b227_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b227_c0 : nS_st7_b227_c1;
  assign nS_st8_b228_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b228_c0 : nS_st7_b228_c1;
  assign nS_st8_b229_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b229_c0 : nS_st7_b229_c1;
  assign nS_st8_b230_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b230_c0 : nS_st7_b230_c1;
  assign nS_st8_b231_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b231_c0 : nS_st7_b231_c1;
  assign nS_st8_b232_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b232_c0 : nS_st7_b232_c1;
  assign nS_st8_b233_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b233_c0 : nS_st7_b233_c1;
  assign nS_st8_b234_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b234_c0 : nS_st7_b234_c1;
  assign nS_st8_b235_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b235_c0 : nS_st7_b235_c1;
  assign nS_st8_b236_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b236_c0 : nS_st7_b236_c1;
  assign nS_st8_b237_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b237_c0 : nS_st7_b237_c1;
  assign nS_st8_b238_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b238_c0 : nS_st7_b238_c1;
  assign nS_st8_b239_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b239_c0 : nS_st7_b239_c1;
  assign nS_st8_b240_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b240_c0 : nS_st7_b240_c1;
  assign nS_st8_b241_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b241_c0 : nS_st7_b241_c1;
  assign nS_st8_b242_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b242_c0 : nS_st7_b242_c1;
  assign nS_st8_b243_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b243_c0 : nS_st7_b243_c1;
  assign nS_st8_b244_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b244_c0 : nS_st7_b244_c1;
  assign nS_st8_b245_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b245_c0 : nS_st7_b245_c1;
  assign nS_st8_b246_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b246_c0 : nS_st7_b246_c1;
  assign nS_st8_b247_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b247_c0 : nS_st7_b247_c1;
  assign nS_st8_b248_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b248_c0 : nS_st7_b248_c1;
  assign nS_st8_b249_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b249_c0 : nS_st7_b249_c1;
  assign nS_st8_b250_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b250_c0 : nS_st7_b250_c1;
  assign nS_st8_b251_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b251_c0 : nS_st7_b251_c1;
  assign nS_st8_b252_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b252_c0 : nS_st7_b252_c1;
  assign nS_st8_b253_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b253_c0 : nS_st7_b253_c1;
  assign nS_st8_b254_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b254_c0 : nS_st7_b254_c1;
  assign nS_st8_b255_c0 = (nC_st7_b191_c0 == 0) ? nS_st7_b255_c0 : nS_st7_b255_c1;
  assign nS_st8_b0_c1 = nS_st7_b0_c1;
  assign nS_st8_b1_c1 = nS_st7_b1_c1;
  assign nS_st8_b2_c1 = nS_st7_b2_c1;
  assign nS_st8_b3_c1 = nS_st7_b3_c1;
  assign nS_st8_b4_c1 = nS_st7_b4_c1;
  assign nS_st8_b5_c1 = nS_st7_b5_c1;
  assign nS_st8_b6_c1 = nS_st7_b6_c1;
  assign nS_st8_b7_c1 = nS_st7_b7_c1;
  assign nS_st8_b8_c1 = nS_st7_b8_c1;
  assign nS_st8_b9_c1 = nS_st7_b9_c1;
  assign nS_st8_b10_c1 = nS_st7_b10_c1;
  assign nS_st8_b11_c1 = nS_st7_b11_c1;
  assign nS_st8_b12_c1 = nS_st7_b12_c1;
  assign nS_st8_b13_c1 = nS_st7_b13_c1;
  assign nS_st8_b14_c1 = nS_st7_b14_c1;
  assign nS_st8_b15_c1 = nS_st7_b15_c1;
  assign nS_st8_b16_c1 = nS_st7_b16_c1;
  assign nS_st8_b17_c1 = nS_st7_b17_c1;
  assign nS_st8_b18_c1 = nS_st7_b18_c1;
  assign nS_st8_b19_c1 = nS_st7_b19_c1;
  assign nS_st8_b20_c1 = nS_st7_b20_c1;
  assign nS_st8_b21_c1 = nS_st7_b21_c1;
  assign nS_st8_b22_c1 = nS_st7_b22_c1;
  assign nS_st8_b23_c1 = nS_st7_b23_c1;
  assign nS_st8_b24_c1 = nS_st7_b24_c1;
  assign nS_st8_b25_c1 = nS_st7_b25_c1;
  assign nS_st8_b26_c1 = nS_st7_b26_c1;
  assign nS_st8_b27_c1 = nS_st7_b27_c1;
  assign nS_st8_b28_c1 = nS_st7_b28_c1;
  assign nS_st8_b29_c1 = nS_st7_b29_c1;
  assign nS_st8_b30_c1 = nS_st7_b30_c1;
  assign nS_st8_b31_c1 = nS_st7_b31_c1;
  assign nS_st8_b32_c1 = nS_st7_b32_c1;
  assign nS_st8_b33_c1 = nS_st7_b33_c1;
  assign nS_st8_b34_c1 = nS_st7_b34_c1;
  assign nS_st8_b35_c1 = nS_st7_b35_c1;
  assign nS_st8_b36_c1 = nS_st7_b36_c1;
  assign nS_st8_b37_c1 = nS_st7_b37_c1;
  assign nS_st8_b38_c1 = nS_st7_b38_c1;
  assign nS_st8_b39_c1 = nS_st7_b39_c1;
  assign nS_st8_b40_c1 = nS_st7_b40_c1;
  assign nS_st8_b41_c1 = nS_st7_b41_c1;
  assign nS_st8_b42_c1 = nS_st7_b42_c1;
  assign nS_st8_b43_c1 = nS_st7_b43_c1;
  assign nS_st8_b44_c1 = nS_st7_b44_c1;
  assign nS_st8_b45_c1 = nS_st7_b45_c1;
  assign nS_st8_b46_c1 = nS_st7_b46_c1;
  assign nS_st8_b47_c1 = nS_st7_b47_c1;
  assign nS_st8_b48_c1 = nS_st7_b48_c1;
  assign nS_st8_b49_c1 = nS_st7_b49_c1;
  assign nS_st8_b50_c1 = nS_st7_b50_c1;
  assign nS_st8_b51_c1 = nS_st7_b51_c1;
  assign nS_st8_b52_c1 = nS_st7_b52_c1;
  assign nS_st8_b53_c1 = nS_st7_b53_c1;
  assign nS_st8_b54_c1 = nS_st7_b54_c1;
  assign nS_st8_b55_c1 = nS_st7_b55_c1;
  assign nS_st8_b56_c1 = nS_st7_b56_c1;
  assign nS_st8_b57_c1 = nS_st7_b57_c1;
  assign nS_st8_b58_c1 = nS_st7_b58_c1;
  assign nS_st8_b59_c1 = nS_st7_b59_c1;
  assign nS_st8_b60_c1 = nS_st7_b60_c1;
  assign nS_st8_b61_c1 = nS_st7_b61_c1;
  assign nS_st8_b62_c1 = nS_st7_b62_c1;
  assign nS_st8_b63_c1 = nS_st7_b63_c1;
  assign nS_st8_b64_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b64_c0 : nS_st7_b64_c1;
  assign nS_st8_b65_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b65_c0 : nS_st7_b65_c1;
  assign nS_st8_b66_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b66_c0 : nS_st7_b66_c1;
  assign nS_st8_b67_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b67_c0 : nS_st7_b67_c1;
  assign nS_st8_b68_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b68_c0 : nS_st7_b68_c1;
  assign nS_st8_b69_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b69_c0 : nS_st7_b69_c1;
  assign nS_st8_b70_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b70_c0 : nS_st7_b70_c1;
  assign nS_st8_b71_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b71_c0 : nS_st7_b71_c1;
  assign nS_st8_b72_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b72_c0 : nS_st7_b72_c1;
  assign nS_st8_b73_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b73_c0 : nS_st7_b73_c1;
  assign nS_st8_b74_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b74_c0 : nS_st7_b74_c1;
  assign nS_st8_b75_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b75_c0 : nS_st7_b75_c1;
  assign nS_st8_b76_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b76_c0 : nS_st7_b76_c1;
  assign nS_st8_b77_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b77_c0 : nS_st7_b77_c1;
  assign nS_st8_b78_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b78_c0 : nS_st7_b78_c1;
  assign nS_st8_b79_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b79_c0 : nS_st7_b79_c1;
  assign nS_st8_b80_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b80_c0 : nS_st7_b80_c1;
  assign nS_st8_b81_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b81_c0 : nS_st7_b81_c1;
  assign nS_st8_b82_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b82_c0 : nS_st7_b82_c1;
  assign nS_st8_b83_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b83_c0 : nS_st7_b83_c1;
  assign nS_st8_b84_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b84_c0 : nS_st7_b84_c1;
  assign nS_st8_b85_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b85_c0 : nS_st7_b85_c1;
  assign nS_st8_b86_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b86_c0 : nS_st7_b86_c1;
  assign nS_st8_b87_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b87_c0 : nS_st7_b87_c1;
  assign nS_st8_b88_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b88_c0 : nS_st7_b88_c1;
  assign nS_st8_b89_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b89_c0 : nS_st7_b89_c1;
  assign nS_st8_b90_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b90_c0 : nS_st7_b90_c1;
  assign nS_st8_b91_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b91_c0 : nS_st7_b91_c1;
  assign nS_st8_b92_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b92_c0 : nS_st7_b92_c1;
  assign nS_st8_b93_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b93_c0 : nS_st7_b93_c1;
  assign nS_st8_b94_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b94_c0 : nS_st7_b94_c1;
  assign nS_st8_b95_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b95_c0 : nS_st7_b95_c1;
  assign nS_st8_b96_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b96_c0 : nS_st7_b96_c1;
  assign nS_st8_b97_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b97_c0 : nS_st7_b97_c1;
  assign nS_st8_b98_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b98_c0 : nS_st7_b98_c1;
  assign nS_st8_b99_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b99_c0 : nS_st7_b99_c1;
  assign nS_st8_b100_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b100_c0 : nS_st7_b100_c1;
  assign nS_st8_b101_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b101_c0 : nS_st7_b101_c1;
  assign nS_st8_b102_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b102_c0 : nS_st7_b102_c1;
  assign nS_st8_b103_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b103_c0 : nS_st7_b103_c1;
  assign nS_st8_b104_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b104_c0 : nS_st7_b104_c1;
  assign nS_st8_b105_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b105_c0 : nS_st7_b105_c1;
  assign nS_st8_b106_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b106_c0 : nS_st7_b106_c1;
  assign nS_st8_b107_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b107_c0 : nS_st7_b107_c1;
  assign nS_st8_b108_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b108_c0 : nS_st7_b108_c1;
  assign nS_st8_b109_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b109_c0 : nS_st7_b109_c1;
  assign nS_st8_b110_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b110_c0 : nS_st7_b110_c1;
  assign nS_st8_b111_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b111_c0 : nS_st7_b111_c1;
  assign nS_st8_b112_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b112_c0 : nS_st7_b112_c1;
  assign nS_st8_b113_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b113_c0 : nS_st7_b113_c1;
  assign nS_st8_b114_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b114_c0 : nS_st7_b114_c1;
  assign nS_st8_b115_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b115_c0 : nS_st7_b115_c1;
  assign nS_st8_b116_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b116_c0 : nS_st7_b116_c1;
  assign nS_st8_b117_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b117_c0 : nS_st7_b117_c1;
  assign nS_st8_b118_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b118_c0 : nS_st7_b118_c1;
  assign nS_st8_b119_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b119_c0 : nS_st7_b119_c1;
  assign nS_st8_b120_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b120_c0 : nS_st7_b120_c1;
  assign nS_st8_b121_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b121_c0 : nS_st7_b121_c1;
  assign nS_st8_b122_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b122_c0 : nS_st7_b122_c1;
  assign nS_st8_b123_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b123_c0 : nS_st7_b123_c1;
  assign nS_st8_b124_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b124_c0 : nS_st7_b124_c1;
  assign nS_st8_b125_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b125_c0 : nS_st7_b125_c1;
  assign nS_st8_b126_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b126_c0 : nS_st7_b126_c1;
  assign nS_st8_b127_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b127_c0 : nS_st7_b127_c1;
  assign nS_st8_b128_c1 = nS_st7_b128_c1;
  assign nS_st8_b129_c1 = nS_st7_b129_c1;
  assign nS_st8_b130_c1 = nS_st7_b130_c1;
  assign nS_st8_b131_c1 = nS_st7_b131_c1;
  assign nS_st8_b132_c1 = nS_st7_b132_c1;
  assign nS_st8_b133_c1 = nS_st7_b133_c1;
  assign nS_st8_b134_c1 = nS_st7_b134_c1;
  assign nS_st8_b135_c1 = nS_st7_b135_c1;
  assign nS_st8_b136_c1 = nS_st7_b136_c1;
  assign nS_st8_b137_c1 = nS_st7_b137_c1;
  assign nS_st8_b138_c1 = nS_st7_b138_c1;
  assign nS_st8_b139_c1 = nS_st7_b139_c1;
  assign nS_st8_b140_c1 = nS_st7_b140_c1;
  assign nS_st8_b141_c1 = nS_st7_b141_c1;
  assign nS_st8_b142_c1 = nS_st7_b142_c1;
  assign nS_st8_b143_c1 = nS_st7_b143_c1;
  assign nS_st8_b144_c1 = nS_st7_b144_c1;
  assign nS_st8_b145_c1 = nS_st7_b145_c1;
  assign nS_st8_b146_c1 = nS_st7_b146_c1;
  assign nS_st8_b147_c1 = nS_st7_b147_c1;
  assign nS_st8_b148_c1 = nS_st7_b148_c1;
  assign nS_st8_b149_c1 = nS_st7_b149_c1;
  assign nS_st8_b150_c1 = nS_st7_b150_c1;
  assign nS_st8_b151_c1 = nS_st7_b151_c1;
  assign nS_st8_b152_c1 = nS_st7_b152_c1;
  assign nS_st8_b153_c1 = nS_st7_b153_c1;
  assign nS_st8_b154_c1 = nS_st7_b154_c1;
  assign nS_st8_b155_c1 = nS_st7_b155_c1;
  assign nS_st8_b156_c1 = nS_st7_b156_c1;
  assign nS_st8_b157_c1 = nS_st7_b157_c1;
  assign nS_st8_b158_c1 = nS_st7_b158_c1;
  assign nS_st8_b159_c1 = nS_st7_b159_c1;
  assign nS_st8_b160_c1 = nS_st7_b160_c1;
  assign nS_st8_b161_c1 = nS_st7_b161_c1;
  assign nS_st8_b162_c1 = nS_st7_b162_c1;
  assign nS_st8_b163_c1 = nS_st7_b163_c1;
  assign nS_st8_b164_c1 = nS_st7_b164_c1;
  assign nS_st8_b165_c1 = nS_st7_b165_c1;
  assign nS_st8_b166_c1 = nS_st7_b166_c1;
  assign nS_st8_b167_c1 = nS_st7_b167_c1;
  assign nS_st8_b168_c1 = nS_st7_b168_c1;
  assign nS_st8_b169_c1 = nS_st7_b169_c1;
  assign nS_st8_b170_c1 = nS_st7_b170_c1;
  assign nS_st8_b171_c1 = nS_st7_b171_c1;
  assign nS_st8_b172_c1 = nS_st7_b172_c1;
  assign nS_st8_b173_c1 = nS_st7_b173_c1;
  assign nS_st8_b174_c1 = nS_st7_b174_c1;
  assign nS_st8_b175_c1 = nS_st7_b175_c1;
  assign nS_st8_b176_c1 = nS_st7_b176_c1;
  assign nS_st8_b177_c1 = nS_st7_b177_c1;
  assign nS_st8_b178_c1 = nS_st7_b178_c1;
  assign nS_st8_b179_c1 = nS_st7_b179_c1;
  assign nS_st8_b180_c1 = nS_st7_b180_c1;
  assign nS_st8_b181_c1 = nS_st7_b181_c1;
  assign nS_st8_b182_c1 = nS_st7_b182_c1;
  assign nS_st8_b183_c1 = nS_st7_b183_c1;
  assign nS_st8_b184_c1 = nS_st7_b184_c1;
  assign nS_st8_b185_c1 = nS_st7_b185_c1;
  assign nS_st8_b186_c1 = nS_st7_b186_c1;
  assign nS_st8_b187_c1 = nS_st7_b187_c1;
  assign nS_st8_b188_c1 = nS_st7_b188_c1;
  assign nS_st8_b189_c1 = nS_st7_b189_c1;
  assign nS_st8_b190_c1 = nS_st7_b190_c1;
  assign nS_st8_b191_c1 = nS_st7_b191_c1;
  assign nS_st8_b192_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b192_c0 : nS_st7_b192_c1;
  assign nS_st8_b193_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b193_c0 : nS_st7_b193_c1;
  assign nS_st8_b194_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b194_c0 : nS_st7_b194_c1;
  assign nS_st8_b195_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b195_c0 : nS_st7_b195_c1;
  assign nS_st8_b196_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b196_c0 : nS_st7_b196_c1;
  assign nS_st8_b197_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b197_c0 : nS_st7_b197_c1;
  assign nS_st8_b198_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b198_c0 : nS_st7_b198_c1;
  assign nS_st8_b199_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b199_c0 : nS_st7_b199_c1;
  assign nS_st8_b200_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b200_c0 : nS_st7_b200_c1;
  assign nS_st8_b201_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b201_c0 : nS_st7_b201_c1;
  assign nS_st8_b202_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b202_c0 : nS_st7_b202_c1;
  assign nS_st8_b203_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b203_c0 : nS_st7_b203_c1;
  assign nS_st8_b204_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b204_c0 : nS_st7_b204_c1;
  assign nS_st8_b205_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b205_c0 : nS_st7_b205_c1;
  assign nS_st8_b206_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b206_c0 : nS_st7_b206_c1;
  assign nS_st8_b207_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b207_c0 : nS_st7_b207_c1;
  assign nS_st8_b208_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b208_c0 : nS_st7_b208_c1;
  assign nS_st8_b209_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b209_c0 : nS_st7_b209_c1;
  assign nS_st8_b210_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b210_c0 : nS_st7_b210_c1;
  assign nS_st8_b211_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b211_c0 : nS_st7_b211_c1;
  assign nS_st8_b212_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b212_c0 : nS_st7_b212_c1;
  assign nS_st8_b213_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b213_c0 : nS_st7_b213_c1;
  assign nS_st8_b214_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b214_c0 : nS_st7_b214_c1;
  assign nS_st8_b215_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b215_c0 : nS_st7_b215_c1;
  assign nS_st8_b216_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b216_c0 : nS_st7_b216_c1;
  assign nS_st8_b217_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b217_c0 : nS_st7_b217_c1;
  assign nS_st8_b218_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b218_c0 : nS_st7_b218_c1;
  assign nS_st8_b219_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b219_c0 : nS_st7_b219_c1;
  assign nS_st8_b220_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b220_c0 : nS_st7_b220_c1;
  assign nS_st8_b221_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b221_c0 : nS_st7_b221_c1;
  assign nS_st8_b222_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b222_c0 : nS_st7_b222_c1;
  assign nS_st8_b223_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b223_c0 : nS_st7_b223_c1;
  assign nS_st8_b224_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b224_c0 : nS_st7_b224_c1;
  assign nS_st8_b225_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b225_c0 : nS_st7_b225_c1;
  assign nS_st8_b226_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b226_c0 : nS_st7_b226_c1;
  assign nS_st8_b227_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b227_c0 : nS_st7_b227_c1;
  assign nS_st8_b228_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b228_c0 : nS_st7_b228_c1;
  assign nS_st8_b229_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b229_c0 : nS_st7_b229_c1;
  assign nS_st8_b230_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b230_c0 : nS_st7_b230_c1;
  assign nS_st8_b231_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b231_c0 : nS_st7_b231_c1;
  assign nS_st8_b232_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b232_c0 : nS_st7_b232_c1;
  assign nS_st8_b233_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b233_c0 : nS_st7_b233_c1;
  assign nS_st8_b234_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b234_c0 : nS_st7_b234_c1;
  assign nS_st8_b235_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b235_c0 : nS_st7_b235_c1;
  assign nS_st8_b236_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b236_c0 : nS_st7_b236_c1;
  assign nS_st8_b237_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b237_c0 : nS_st7_b237_c1;
  assign nS_st8_b238_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b238_c0 : nS_st7_b238_c1;
  assign nS_st8_b239_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b239_c0 : nS_st7_b239_c1;
  assign nS_st8_b240_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b240_c0 : nS_st7_b240_c1;
  assign nS_st8_b241_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b241_c0 : nS_st7_b241_c1;
  assign nS_st8_b242_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b242_c0 : nS_st7_b242_c1;
  assign nS_st8_b243_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b243_c0 : nS_st7_b243_c1;
  assign nS_st8_b244_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b244_c0 : nS_st7_b244_c1;
  assign nS_st8_b245_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b245_c0 : nS_st7_b245_c1;
  assign nS_st8_b246_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b246_c0 : nS_st7_b246_c1;
  assign nS_st8_b247_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b247_c0 : nS_st7_b247_c1;
  assign nS_st8_b248_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b248_c0 : nS_st7_b248_c1;
  assign nS_st8_b249_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b249_c0 : nS_st7_b249_c1;
  assign nS_st8_b250_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b250_c0 : nS_st7_b250_c1;
  assign nS_st8_b251_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b251_c0 : nS_st7_b251_c1;
  assign nS_st8_b252_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b252_c0 : nS_st7_b252_c1;
  assign nS_st8_b253_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b253_c0 : nS_st7_b253_c1;
  assign nS_st8_b254_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b254_c0 : nS_st7_b254_c1;
  assign nS_st8_b255_c1 = (nC_st7_b191_c1 == 0) ? nS_st7_b255_c0 : nS_st7_b255_c1;
  assign nC_st8_b127_c0 = (nC_st7_b63_c0 == 0) ? nC_st7_b127_c0 : nC_st7_b127_c1;
  assign nC_st8_b255_c0 = (nC_st7_b191_c0 == 0) ? nC_st7_b255_c0 : nC_st7_b255_c1;
  assign nC_st8_b127_c1 = (nC_st7_b63_c1 == 0) ? nC_st7_b127_c0 : nC_st7_b127_c1;
  assign nC_st8_b255_c1 = (nC_st7_b191_c1 == 0) ? nC_st7_b255_c0 : nC_st7_b255_c1;

  assign nS_st9_b0_c0 = nS_st8_b0_c0;
  assign nS_st9_b1_c0 = nS_st8_b1_c0;
  assign nS_st9_b2_c0 = nS_st8_b2_c0;
  assign nS_st9_b3_c0 = nS_st8_b3_c0;
  assign nS_st9_b4_c0 = nS_st8_b4_c0;
  assign nS_st9_b5_c0 = nS_st8_b5_c0;
  assign nS_st9_b6_c0 = nS_st8_b6_c0;
  assign nS_st9_b7_c0 = nS_st8_b7_c0;
  assign nS_st9_b8_c0 = nS_st8_b8_c0;
  assign nS_st9_b9_c0 = nS_st8_b9_c0;
  assign nS_st9_b10_c0 = nS_st8_b10_c0;
  assign nS_st9_b11_c0 = nS_st8_b11_c0;
  assign nS_st9_b12_c0 = nS_st8_b12_c0;
  assign nS_st9_b13_c0 = nS_st8_b13_c0;
  assign nS_st9_b14_c0 = nS_st8_b14_c0;
  assign nS_st9_b15_c0 = nS_st8_b15_c0;
  assign nS_st9_b16_c0 = nS_st8_b16_c0;
  assign nS_st9_b17_c0 = nS_st8_b17_c0;
  assign nS_st9_b18_c0 = nS_st8_b18_c0;
  assign nS_st9_b19_c0 = nS_st8_b19_c0;
  assign nS_st9_b20_c0 = nS_st8_b20_c0;
  assign nS_st9_b21_c0 = nS_st8_b21_c0;
  assign nS_st9_b22_c0 = nS_st8_b22_c0;
  assign nS_st9_b23_c0 = nS_st8_b23_c0;
  assign nS_st9_b24_c0 = nS_st8_b24_c0;
  assign nS_st9_b25_c0 = nS_st8_b25_c0;
  assign nS_st9_b26_c0 = nS_st8_b26_c0;
  assign nS_st9_b27_c0 = nS_st8_b27_c0;
  assign nS_st9_b28_c0 = nS_st8_b28_c0;
  assign nS_st9_b29_c0 = nS_st8_b29_c0;
  assign nS_st9_b30_c0 = nS_st8_b30_c0;
  assign nS_st9_b31_c0 = nS_st8_b31_c0;
  assign nS_st9_b32_c0 = nS_st8_b32_c0;
  assign nS_st9_b33_c0 = nS_st8_b33_c0;
  assign nS_st9_b34_c0 = nS_st8_b34_c0;
  assign nS_st9_b35_c0 = nS_st8_b35_c0;
  assign nS_st9_b36_c0 = nS_st8_b36_c0;
  assign nS_st9_b37_c0 = nS_st8_b37_c0;
  assign nS_st9_b38_c0 = nS_st8_b38_c0;
  assign nS_st9_b39_c0 = nS_st8_b39_c0;
  assign nS_st9_b40_c0 = nS_st8_b40_c0;
  assign nS_st9_b41_c0 = nS_st8_b41_c0;
  assign nS_st9_b42_c0 = nS_st8_b42_c0;
  assign nS_st9_b43_c0 = nS_st8_b43_c0;
  assign nS_st9_b44_c0 = nS_st8_b44_c0;
  assign nS_st9_b45_c0 = nS_st8_b45_c0;
  assign nS_st9_b46_c0 = nS_st8_b46_c0;
  assign nS_st9_b47_c0 = nS_st8_b47_c0;
  assign nS_st9_b48_c0 = nS_st8_b48_c0;
  assign nS_st9_b49_c0 = nS_st8_b49_c0;
  assign nS_st9_b50_c0 = nS_st8_b50_c0;
  assign nS_st9_b51_c0 = nS_st8_b51_c0;
  assign nS_st9_b52_c0 = nS_st8_b52_c0;
  assign nS_st9_b53_c0 = nS_st8_b53_c0;
  assign nS_st9_b54_c0 = nS_st8_b54_c0;
  assign nS_st9_b55_c0 = nS_st8_b55_c0;
  assign nS_st9_b56_c0 = nS_st8_b56_c0;
  assign nS_st9_b57_c0 = nS_st8_b57_c0;
  assign nS_st9_b58_c0 = nS_st8_b58_c0;
  assign nS_st9_b59_c0 = nS_st8_b59_c0;
  assign nS_st9_b60_c0 = nS_st8_b60_c0;
  assign nS_st9_b61_c0 = nS_st8_b61_c0;
  assign nS_st9_b62_c0 = nS_st8_b62_c0;
  assign nS_st9_b63_c0 = nS_st8_b63_c0;
  assign nS_st9_b64_c0 = nS_st8_b64_c0;
  assign nS_st9_b65_c0 = nS_st8_b65_c0;
  assign nS_st9_b66_c0 = nS_st8_b66_c0;
  assign nS_st9_b67_c0 = nS_st8_b67_c0;
  assign nS_st9_b68_c0 = nS_st8_b68_c0;
  assign nS_st9_b69_c0 = nS_st8_b69_c0;
  assign nS_st9_b70_c0 = nS_st8_b70_c0;
  assign nS_st9_b71_c0 = nS_st8_b71_c0;
  assign nS_st9_b72_c0 = nS_st8_b72_c0;
  assign nS_st9_b73_c0 = nS_st8_b73_c0;
  assign nS_st9_b74_c0 = nS_st8_b74_c0;
  assign nS_st9_b75_c0 = nS_st8_b75_c0;
  assign nS_st9_b76_c0 = nS_st8_b76_c0;
  assign nS_st9_b77_c0 = nS_st8_b77_c0;
  assign nS_st9_b78_c0 = nS_st8_b78_c0;
  assign nS_st9_b79_c0 = nS_st8_b79_c0;
  assign nS_st9_b80_c0 = nS_st8_b80_c0;
  assign nS_st9_b81_c0 = nS_st8_b81_c0;
  assign nS_st9_b82_c0 = nS_st8_b82_c0;
  assign nS_st9_b83_c0 = nS_st8_b83_c0;
  assign nS_st9_b84_c0 = nS_st8_b84_c0;
  assign nS_st9_b85_c0 = nS_st8_b85_c0;
  assign nS_st9_b86_c0 = nS_st8_b86_c0;
  assign nS_st9_b87_c0 = nS_st8_b87_c0;
  assign nS_st9_b88_c0 = nS_st8_b88_c0;
  assign nS_st9_b89_c0 = nS_st8_b89_c0;
  assign nS_st9_b90_c0 = nS_st8_b90_c0;
  assign nS_st9_b91_c0 = nS_st8_b91_c0;
  assign nS_st9_b92_c0 = nS_st8_b92_c0;
  assign nS_st9_b93_c0 = nS_st8_b93_c0;
  assign nS_st9_b94_c0 = nS_st8_b94_c0;
  assign nS_st9_b95_c0 = nS_st8_b95_c0;
  assign nS_st9_b96_c0 = nS_st8_b96_c0;
  assign nS_st9_b97_c0 = nS_st8_b97_c0;
  assign nS_st9_b98_c0 = nS_st8_b98_c0;
  assign nS_st9_b99_c0 = nS_st8_b99_c0;
  assign nS_st9_b100_c0 = nS_st8_b100_c0;
  assign nS_st9_b101_c0 = nS_st8_b101_c0;
  assign nS_st9_b102_c0 = nS_st8_b102_c0;
  assign nS_st9_b103_c0 = nS_st8_b103_c0;
  assign nS_st9_b104_c0 = nS_st8_b104_c0;
  assign nS_st9_b105_c0 = nS_st8_b105_c0;
  assign nS_st9_b106_c0 = nS_st8_b106_c0;
  assign nS_st9_b107_c0 = nS_st8_b107_c0;
  assign nS_st9_b108_c0 = nS_st8_b108_c0;
  assign nS_st9_b109_c0 = nS_st8_b109_c0;
  assign nS_st9_b110_c0 = nS_st8_b110_c0;
  assign nS_st9_b111_c0 = nS_st8_b111_c0;
  assign nS_st9_b112_c0 = nS_st8_b112_c0;
  assign nS_st9_b113_c0 = nS_st8_b113_c0;
  assign nS_st9_b114_c0 = nS_st8_b114_c0;
  assign nS_st9_b115_c0 = nS_st8_b115_c0;
  assign nS_st9_b116_c0 = nS_st8_b116_c0;
  assign nS_st9_b117_c0 = nS_st8_b117_c0;
  assign nS_st9_b118_c0 = nS_st8_b118_c0;
  assign nS_st9_b119_c0 = nS_st8_b119_c0;
  assign nS_st9_b120_c0 = nS_st8_b120_c0;
  assign nS_st9_b121_c0 = nS_st8_b121_c0;
  assign nS_st9_b122_c0 = nS_st8_b122_c0;
  assign nS_st9_b123_c0 = nS_st8_b123_c0;
  assign nS_st9_b124_c0 = nS_st8_b124_c0;
  assign nS_st9_b125_c0 = nS_st8_b125_c0;
  assign nS_st9_b126_c0 = nS_st8_b126_c0;
  assign nS_st9_b127_c0 = nS_st8_b127_c0;
  assign nS_st9_b128_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b128_c0 : nS_st8_b128_c1;
  assign nS_st9_b129_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b129_c0 : nS_st8_b129_c1;
  assign nS_st9_b130_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b130_c0 : nS_st8_b130_c1;
  assign nS_st9_b131_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b131_c0 : nS_st8_b131_c1;
  assign nS_st9_b132_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b132_c0 : nS_st8_b132_c1;
  assign nS_st9_b133_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b133_c0 : nS_st8_b133_c1;
  assign nS_st9_b134_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b134_c0 : nS_st8_b134_c1;
  assign nS_st9_b135_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b135_c0 : nS_st8_b135_c1;
  assign nS_st9_b136_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b136_c0 : nS_st8_b136_c1;
  assign nS_st9_b137_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b137_c0 : nS_st8_b137_c1;
  assign nS_st9_b138_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b138_c0 : nS_st8_b138_c1;
  assign nS_st9_b139_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b139_c0 : nS_st8_b139_c1;
  assign nS_st9_b140_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b140_c0 : nS_st8_b140_c1;
  assign nS_st9_b141_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b141_c0 : nS_st8_b141_c1;
  assign nS_st9_b142_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b142_c0 : nS_st8_b142_c1;
  assign nS_st9_b143_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b143_c0 : nS_st8_b143_c1;
  assign nS_st9_b144_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b144_c0 : nS_st8_b144_c1;
  assign nS_st9_b145_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b145_c0 : nS_st8_b145_c1;
  assign nS_st9_b146_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b146_c0 : nS_st8_b146_c1;
  assign nS_st9_b147_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b147_c0 : nS_st8_b147_c1;
  assign nS_st9_b148_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b148_c0 : nS_st8_b148_c1;
  assign nS_st9_b149_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b149_c0 : nS_st8_b149_c1;
  assign nS_st9_b150_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b150_c0 : nS_st8_b150_c1;
  assign nS_st9_b151_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b151_c0 : nS_st8_b151_c1;
  assign nS_st9_b152_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b152_c0 : nS_st8_b152_c1;
  assign nS_st9_b153_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b153_c0 : nS_st8_b153_c1;
  assign nS_st9_b154_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b154_c0 : nS_st8_b154_c1;
  assign nS_st9_b155_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b155_c0 : nS_st8_b155_c1;
  assign nS_st9_b156_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b156_c0 : nS_st8_b156_c1;
  assign nS_st9_b157_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b157_c0 : nS_st8_b157_c1;
  assign nS_st9_b158_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b158_c0 : nS_st8_b158_c1;
  assign nS_st9_b159_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b159_c0 : nS_st8_b159_c1;
  assign nS_st9_b160_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b160_c0 : nS_st8_b160_c1;
  assign nS_st9_b161_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b161_c0 : nS_st8_b161_c1;
  assign nS_st9_b162_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b162_c0 : nS_st8_b162_c1;
  assign nS_st9_b163_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b163_c0 : nS_st8_b163_c1;
  assign nS_st9_b164_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b164_c0 : nS_st8_b164_c1;
  assign nS_st9_b165_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b165_c0 : nS_st8_b165_c1;
  assign nS_st9_b166_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b166_c0 : nS_st8_b166_c1;
  assign nS_st9_b167_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b167_c0 : nS_st8_b167_c1;
  assign nS_st9_b168_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b168_c0 : nS_st8_b168_c1;
  assign nS_st9_b169_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b169_c0 : nS_st8_b169_c1;
  assign nS_st9_b170_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b170_c0 : nS_st8_b170_c1;
  assign nS_st9_b171_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b171_c0 : nS_st8_b171_c1;
  assign nS_st9_b172_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b172_c0 : nS_st8_b172_c1;
  assign nS_st9_b173_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b173_c0 : nS_st8_b173_c1;
  assign nS_st9_b174_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b174_c0 : nS_st8_b174_c1;
  assign nS_st9_b175_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b175_c0 : nS_st8_b175_c1;
  assign nS_st9_b176_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b176_c0 : nS_st8_b176_c1;
  assign nS_st9_b177_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b177_c0 : nS_st8_b177_c1;
  assign nS_st9_b178_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b178_c0 : nS_st8_b178_c1;
  assign nS_st9_b179_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b179_c0 : nS_st8_b179_c1;
  assign nS_st9_b180_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b180_c0 : nS_st8_b180_c1;
  assign nS_st9_b181_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b181_c0 : nS_st8_b181_c1;
  assign nS_st9_b182_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b182_c0 : nS_st8_b182_c1;
  assign nS_st9_b183_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b183_c0 : nS_st8_b183_c1;
  assign nS_st9_b184_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b184_c0 : nS_st8_b184_c1;
  assign nS_st9_b185_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b185_c0 : nS_st8_b185_c1;
  assign nS_st9_b186_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b186_c0 : nS_st8_b186_c1;
  assign nS_st9_b187_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b187_c0 : nS_st8_b187_c1;
  assign nS_st9_b188_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b188_c0 : nS_st8_b188_c1;
  assign nS_st9_b189_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b189_c0 : nS_st8_b189_c1;
  assign nS_st9_b190_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b190_c0 : nS_st8_b190_c1;
  assign nS_st9_b191_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b191_c0 : nS_st8_b191_c1;
  assign nS_st9_b192_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b192_c0 : nS_st8_b192_c1;
  assign nS_st9_b193_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b193_c0 : nS_st8_b193_c1;
  assign nS_st9_b194_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b194_c0 : nS_st8_b194_c1;
  assign nS_st9_b195_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b195_c0 : nS_st8_b195_c1;
  assign nS_st9_b196_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b196_c0 : nS_st8_b196_c1;
  assign nS_st9_b197_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b197_c0 : nS_st8_b197_c1;
  assign nS_st9_b198_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b198_c0 : nS_st8_b198_c1;
  assign nS_st9_b199_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b199_c0 : nS_st8_b199_c1;
  assign nS_st9_b200_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b200_c0 : nS_st8_b200_c1;
  assign nS_st9_b201_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b201_c0 : nS_st8_b201_c1;
  assign nS_st9_b202_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b202_c0 : nS_st8_b202_c1;
  assign nS_st9_b203_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b203_c0 : nS_st8_b203_c1;
  assign nS_st9_b204_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b204_c0 : nS_st8_b204_c1;
  assign nS_st9_b205_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b205_c0 : nS_st8_b205_c1;
  assign nS_st9_b206_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b206_c0 : nS_st8_b206_c1;
  assign nS_st9_b207_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b207_c0 : nS_st8_b207_c1;
  assign nS_st9_b208_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b208_c0 : nS_st8_b208_c1;
  assign nS_st9_b209_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b209_c0 : nS_st8_b209_c1;
  assign nS_st9_b210_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b210_c0 : nS_st8_b210_c1;
  assign nS_st9_b211_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b211_c0 : nS_st8_b211_c1;
  assign nS_st9_b212_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b212_c0 : nS_st8_b212_c1;
  assign nS_st9_b213_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b213_c0 : nS_st8_b213_c1;
  assign nS_st9_b214_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b214_c0 : nS_st8_b214_c1;
  assign nS_st9_b215_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b215_c0 : nS_st8_b215_c1;
  assign nS_st9_b216_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b216_c0 : nS_st8_b216_c1;
  assign nS_st9_b217_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b217_c0 : nS_st8_b217_c1;
  assign nS_st9_b218_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b218_c0 : nS_st8_b218_c1;
  assign nS_st9_b219_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b219_c0 : nS_st8_b219_c1;
  assign nS_st9_b220_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b220_c0 : nS_st8_b220_c1;
  assign nS_st9_b221_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b221_c0 : nS_st8_b221_c1;
  assign nS_st9_b222_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b222_c0 : nS_st8_b222_c1;
  assign nS_st9_b223_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b223_c0 : nS_st8_b223_c1;
  assign nS_st9_b224_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b224_c0 : nS_st8_b224_c1;
  assign nS_st9_b225_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b225_c0 : nS_st8_b225_c1;
  assign nS_st9_b226_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b226_c0 : nS_st8_b226_c1;
  assign nS_st9_b227_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b227_c0 : nS_st8_b227_c1;
  assign nS_st9_b228_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b228_c0 : nS_st8_b228_c1;
  assign nS_st9_b229_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b229_c0 : nS_st8_b229_c1;
  assign nS_st9_b230_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b230_c0 : nS_st8_b230_c1;
  assign nS_st9_b231_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b231_c0 : nS_st8_b231_c1;
  assign nS_st9_b232_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b232_c0 : nS_st8_b232_c1;
  assign nS_st9_b233_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b233_c0 : nS_st8_b233_c1;
  assign nS_st9_b234_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b234_c0 : nS_st8_b234_c1;
  assign nS_st9_b235_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b235_c0 : nS_st8_b235_c1;
  assign nS_st9_b236_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b236_c0 : nS_st8_b236_c1;
  assign nS_st9_b237_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b237_c0 : nS_st8_b237_c1;
  assign nS_st9_b238_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b238_c0 : nS_st8_b238_c1;
  assign nS_st9_b239_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b239_c0 : nS_st8_b239_c1;
  assign nS_st9_b240_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b240_c0 : nS_st8_b240_c1;
  assign nS_st9_b241_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b241_c0 : nS_st8_b241_c1;
  assign nS_st9_b242_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b242_c0 : nS_st8_b242_c1;
  assign nS_st9_b243_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b243_c0 : nS_st8_b243_c1;
  assign nS_st9_b244_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b244_c0 : nS_st8_b244_c1;
  assign nS_st9_b245_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b245_c0 : nS_st8_b245_c1;
  assign nS_st9_b246_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b246_c0 : nS_st8_b246_c1;
  assign nS_st9_b247_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b247_c0 : nS_st8_b247_c1;
  assign nS_st9_b248_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b248_c0 : nS_st8_b248_c1;
  assign nS_st9_b249_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b249_c0 : nS_st8_b249_c1;
  assign nS_st9_b250_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b250_c0 : nS_st8_b250_c1;
  assign nS_st9_b251_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b251_c0 : nS_st8_b251_c1;
  assign nS_st9_b252_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b252_c0 : nS_st8_b252_c1;
  assign nS_st9_b253_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b253_c0 : nS_st8_b253_c1;
  assign nS_st9_b254_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b254_c0 : nS_st8_b254_c1;
  assign nS_st9_b255_c0 = (nC_st8_b127_c0 == 0) ? nS_st8_b255_c0 : nS_st8_b255_c1;
  assign nS_st9_b0_c1 = nS_st8_b0_c1;
  assign nS_st9_b1_c1 = nS_st8_b1_c1;
  assign nS_st9_b2_c1 = nS_st8_b2_c1;
  assign nS_st9_b3_c1 = nS_st8_b3_c1;
  assign nS_st9_b4_c1 = nS_st8_b4_c1;
  assign nS_st9_b5_c1 = nS_st8_b5_c1;
  assign nS_st9_b6_c1 = nS_st8_b6_c1;
  assign nS_st9_b7_c1 = nS_st8_b7_c1;
  assign nS_st9_b8_c1 = nS_st8_b8_c1;
  assign nS_st9_b9_c1 = nS_st8_b9_c1;
  assign nS_st9_b10_c1 = nS_st8_b10_c1;
  assign nS_st9_b11_c1 = nS_st8_b11_c1;
  assign nS_st9_b12_c1 = nS_st8_b12_c1;
  assign nS_st9_b13_c1 = nS_st8_b13_c1;
  assign nS_st9_b14_c1 = nS_st8_b14_c1;
  assign nS_st9_b15_c1 = nS_st8_b15_c1;
  assign nS_st9_b16_c1 = nS_st8_b16_c1;
  assign nS_st9_b17_c1 = nS_st8_b17_c1;
  assign nS_st9_b18_c1 = nS_st8_b18_c1;
  assign nS_st9_b19_c1 = nS_st8_b19_c1;
  assign nS_st9_b20_c1 = nS_st8_b20_c1;
  assign nS_st9_b21_c1 = nS_st8_b21_c1;
  assign nS_st9_b22_c1 = nS_st8_b22_c1;
  assign nS_st9_b23_c1 = nS_st8_b23_c1;
  assign nS_st9_b24_c1 = nS_st8_b24_c1;
  assign nS_st9_b25_c1 = nS_st8_b25_c1;
  assign nS_st9_b26_c1 = nS_st8_b26_c1;
  assign nS_st9_b27_c1 = nS_st8_b27_c1;
  assign nS_st9_b28_c1 = nS_st8_b28_c1;
  assign nS_st9_b29_c1 = nS_st8_b29_c1;
  assign nS_st9_b30_c1 = nS_st8_b30_c1;
  assign nS_st9_b31_c1 = nS_st8_b31_c1;
  assign nS_st9_b32_c1 = nS_st8_b32_c1;
  assign nS_st9_b33_c1 = nS_st8_b33_c1;
  assign nS_st9_b34_c1 = nS_st8_b34_c1;
  assign nS_st9_b35_c1 = nS_st8_b35_c1;
  assign nS_st9_b36_c1 = nS_st8_b36_c1;
  assign nS_st9_b37_c1 = nS_st8_b37_c1;
  assign nS_st9_b38_c1 = nS_st8_b38_c1;
  assign nS_st9_b39_c1 = nS_st8_b39_c1;
  assign nS_st9_b40_c1 = nS_st8_b40_c1;
  assign nS_st9_b41_c1 = nS_st8_b41_c1;
  assign nS_st9_b42_c1 = nS_st8_b42_c1;
  assign nS_st9_b43_c1 = nS_st8_b43_c1;
  assign nS_st9_b44_c1 = nS_st8_b44_c1;
  assign nS_st9_b45_c1 = nS_st8_b45_c1;
  assign nS_st9_b46_c1 = nS_st8_b46_c1;
  assign nS_st9_b47_c1 = nS_st8_b47_c1;
  assign nS_st9_b48_c1 = nS_st8_b48_c1;
  assign nS_st9_b49_c1 = nS_st8_b49_c1;
  assign nS_st9_b50_c1 = nS_st8_b50_c1;
  assign nS_st9_b51_c1 = nS_st8_b51_c1;
  assign nS_st9_b52_c1 = nS_st8_b52_c1;
  assign nS_st9_b53_c1 = nS_st8_b53_c1;
  assign nS_st9_b54_c1 = nS_st8_b54_c1;
  assign nS_st9_b55_c1 = nS_st8_b55_c1;
  assign nS_st9_b56_c1 = nS_st8_b56_c1;
  assign nS_st9_b57_c1 = nS_st8_b57_c1;
  assign nS_st9_b58_c1 = nS_st8_b58_c1;
  assign nS_st9_b59_c1 = nS_st8_b59_c1;
  assign nS_st9_b60_c1 = nS_st8_b60_c1;
  assign nS_st9_b61_c1 = nS_st8_b61_c1;
  assign nS_st9_b62_c1 = nS_st8_b62_c1;
  assign nS_st9_b63_c1 = nS_st8_b63_c1;
  assign nS_st9_b64_c1 = nS_st8_b64_c1;
  assign nS_st9_b65_c1 = nS_st8_b65_c1;
  assign nS_st9_b66_c1 = nS_st8_b66_c1;
  assign nS_st9_b67_c1 = nS_st8_b67_c1;
  assign nS_st9_b68_c1 = nS_st8_b68_c1;
  assign nS_st9_b69_c1 = nS_st8_b69_c1;
  assign nS_st9_b70_c1 = nS_st8_b70_c1;
  assign nS_st9_b71_c1 = nS_st8_b71_c1;
  assign nS_st9_b72_c1 = nS_st8_b72_c1;
  assign nS_st9_b73_c1 = nS_st8_b73_c1;
  assign nS_st9_b74_c1 = nS_st8_b74_c1;
  assign nS_st9_b75_c1 = nS_st8_b75_c1;
  assign nS_st9_b76_c1 = nS_st8_b76_c1;
  assign nS_st9_b77_c1 = nS_st8_b77_c1;
  assign nS_st9_b78_c1 = nS_st8_b78_c1;
  assign nS_st9_b79_c1 = nS_st8_b79_c1;
  assign nS_st9_b80_c1 = nS_st8_b80_c1;
  assign nS_st9_b81_c1 = nS_st8_b81_c1;
  assign nS_st9_b82_c1 = nS_st8_b82_c1;
  assign nS_st9_b83_c1 = nS_st8_b83_c1;
  assign nS_st9_b84_c1 = nS_st8_b84_c1;
  assign nS_st9_b85_c1 = nS_st8_b85_c1;
  assign nS_st9_b86_c1 = nS_st8_b86_c1;
  assign nS_st9_b87_c1 = nS_st8_b87_c1;
  assign nS_st9_b88_c1 = nS_st8_b88_c1;
  assign nS_st9_b89_c1 = nS_st8_b89_c1;
  assign nS_st9_b90_c1 = nS_st8_b90_c1;
  assign nS_st9_b91_c1 = nS_st8_b91_c1;
  assign nS_st9_b92_c1 = nS_st8_b92_c1;
  assign nS_st9_b93_c1 = nS_st8_b93_c1;
  assign nS_st9_b94_c1 = nS_st8_b94_c1;
  assign nS_st9_b95_c1 = nS_st8_b95_c1;
  assign nS_st9_b96_c1 = nS_st8_b96_c1;
  assign nS_st9_b97_c1 = nS_st8_b97_c1;
  assign nS_st9_b98_c1 = nS_st8_b98_c1;
  assign nS_st9_b99_c1 = nS_st8_b99_c1;
  assign nS_st9_b100_c1 = nS_st8_b100_c1;
  assign nS_st9_b101_c1 = nS_st8_b101_c1;
  assign nS_st9_b102_c1 = nS_st8_b102_c1;
  assign nS_st9_b103_c1 = nS_st8_b103_c1;
  assign nS_st9_b104_c1 = nS_st8_b104_c1;
  assign nS_st9_b105_c1 = nS_st8_b105_c1;
  assign nS_st9_b106_c1 = nS_st8_b106_c1;
  assign nS_st9_b107_c1 = nS_st8_b107_c1;
  assign nS_st9_b108_c1 = nS_st8_b108_c1;
  assign nS_st9_b109_c1 = nS_st8_b109_c1;
  assign nS_st9_b110_c1 = nS_st8_b110_c1;
  assign nS_st9_b111_c1 = nS_st8_b111_c1;
  assign nS_st9_b112_c1 = nS_st8_b112_c1;
  assign nS_st9_b113_c1 = nS_st8_b113_c1;
  assign nS_st9_b114_c1 = nS_st8_b114_c1;
  assign nS_st9_b115_c1 = nS_st8_b115_c1;
  assign nS_st9_b116_c1 = nS_st8_b116_c1;
  assign nS_st9_b117_c1 = nS_st8_b117_c1;
  assign nS_st9_b118_c1 = nS_st8_b118_c1;
  assign nS_st9_b119_c1 = nS_st8_b119_c1;
  assign nS_st9_b120_c1 = nS_st8_b120_c1;
  assign nS_st9_b121_c1 = nS_st8_b121_c1;
  assign nS_st9_b122_c1 = nS_st8_b122_c1;
  assign nS_st9_b123_c1 = nS_st8_b123_c1;
  assign nS_st9_b124_c1 = nS_st8_b124_c1;
  assign nS_st9_b125_c1 = nS_st8_b125_c1;
  assign nS_st9_b126_c1 = nS_st8_b126_c1;
  assign nS_st9_b127_c1 = nS_st8_b127_c1;
  assign nS_st9_b128_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b128_c0 : nS_st8_b128_c1;
  assign nS_st9_b129_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b129_c0 : nS_st8_b129_c1;
  assign nS_st9_b130_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b130_c0 : nS_st8_b130_c1;
  assign nS_st9_b131_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b131_c0 : nS_st8_b131_c1;
  assign nS_st9_b132_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b132_c0 : nS_st8_b132_c1;
  assign nS_st9_b133_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b133_c0 : nS_st8_b133_c1;
  assign nS_st9_b134_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b134_c0 : nS_st8_b134_c1;
  assign nS_st9_b135_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b135_c0 : nS_st8_b135_c1;
  assign nS_st9_b136_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b136_c0 : nS_st8_b136_c1;
  assign nS_st9_b137_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b137_c0 : nS_st8_b137_c1;
  assign nS_st9_b138_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b138_c0 : nS_st8_b138_c1;
  assign nS_st9_b139_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b139_c0 : nS_st8_b139_c1;
  assign nS_st9_b140_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b140_c0 : nS_st8_b140_c1;
  assign nS_st9_b141_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b141_c0 : nS_st8_b141_c1;
  assign nS_st9_b142_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b142_c0 : nS_st8_b142_c1;
  assign nS_st9_b143_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b143_c0 : nS_st8_b143_c1;
  assign nS_st9_b144_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b144_c0 : nS_st8_b144_c1;
  assign nS_st9_b145_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b145_c0 : nS_st8_b145_c1;
  assign nS_st9_b146_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b146_c0 : nS_st8_b146_c1;
  assign nS_st9_b147_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b147_c0 : nS_st8_b147_c1;
  assign nS_st9_b148_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b148_c0 : nS_st8_b148_c1;
  assign nS_st9_b149_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b149_c0 : nS_st8_b149_c1;
  assign nS_st9_b150_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b150_c0 : nS_st8_b150_c1;
  assign nS_st9_b151_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b151_c0 : nS_st8_b151_c1;
  assign nS_st9_b152_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b152_c0 : nS_st8_b152_c1;
  assign nS_st9_b153_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b153_c0 : nS_st8_b153_c1;
  assign nS_st9_b154_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b154_c0 : nS_st8_b154_c1;
  assign nS_st9_b155_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b155_c0 : nS_st8_b155_c1;
  assign nS_st9_b156_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b156_c0 : nS_st8_b156_c1;
  assign nS_st9_b157_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b157_c0 : nS_st8_b157_c1;
  assign nS_st9_b158_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b158_c0 : nS_st8_b158_c1;
  assign nS_st9_b159_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b159_c0 : nS_st8_b159_c1;
  assign nS_st9_b160_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b160_c0 : nS_st8_b160_c1;
  assign nS_st9_b161_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b161_c0 : nS_st8_b161_c1;
  assign nS_st9_b162_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b162_c0 : nS_st8_b162_c1;
  assign nS_st9_b163_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b163_c0 : nS_st8_b163_c1;
  assign nS_st9_b164_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b164_c0 : nS_st8_b164_c1;
  assign nS_st9_b165_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b165_c0 : nS_st8_b165_c1;
  assign nS_st9_b166_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b166_c0 : nS_st8_b166_c1;
  assign nS_st9_b167_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b167_c0 : nS_st8_b167_c1;
  assign nS_st9_b168_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b168_c0 : nS_st8_b168_c1;
  assign nS_st9_b169_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b169_c0 : nS_st8_b169_c1;
  assign nS_st9_b170_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b170_c0 : nS_st8_b170_c1;
  assign nS_st9_b171_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b171_c0 : nS_st8_b171_c1;
  assign nS_st9_b172_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b172_c0 : nS_st8_b172_c1;
  assign nS_st9_b173_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b173_c0 : nS_st8_b173_c1;
  assign nS_st9_b174_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b174_c0 : nS_st8_b174_c1;
  assign nS_st9_b175_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b175_c0 : nS_st8_b175_c1;
  assign nS_st9_b176_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b176_c0 : nS_st8_b176_c1;
  assign nS_st9_b177_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b177_c0 : nS_st8_b177_c1;
  assign nS_st9_b178_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b178_c0 : nS_st8_b178_c1;
  assign nS_st9_b179_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b179_c0 : nS_st8_b179_c1;
  assign nS_st9_b180_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b180_c0 : nS_st8_b180_c1;
  assign nS_st9_b181_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b181_c0 : nS_st8_b181_c1;
  assign nS_st9_b182_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b182_c0 : nS_st8_b182_c1;
  assign nS_st9_b183_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b183_c0 : nS_st8_b183_c1;
  assign nS_st9_b184_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b184_c0 : nS_st8_b184_c1;
  assign nS_st9_b185_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b185_c0 : nS_st8_b185_c1;
  assign nS_st9_b186_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b186_c0 : nS_st8_b186_c1;
  assign nS_st9_b187_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b187_c0 : nS_st8_b187_c1;
  assign nS_st9_b188_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b188_c0 : nS_st8_b188_c1;
  assign nS_st9_b189_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b189_c0 : nS_st8_b189_c1;
  assign nS_st9_b190_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b190_c0 : nS_st8_b190_c1;
  assign nS_st9_b191_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b191_c0 : nS_st8_b191_c1;
  assign nS_st9_b192_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b192_c0 : nS_st8_b192_c1;
  assign nS_st9_b193_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b193_c0 : nS_st8_b193_c1;
  assign nS_st9_b194_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b194_c0 : nS_st8_b194_c1;
  assign nS_st9_b195_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b195_c0 : nS_st8_b195_c1;
  assign nS_st9_b196_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b196_c0 : nS_st8_b196_c1;
  assign nS_st9_b197_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b197_c0 : nS_st8_b197_c1;
  assign nS_st9_b198_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b198_c0 : nS_st8_b198_c1;
  assign nS_st9_b199_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b199_c0 : nS_st8_b199_c1;
  assign nS_st9_b200_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b200_c0 : nS_st8_b200_c1;
  assign nS_st9_b201_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b201_c0 : nS_st8_b201_c1;
  assign nS_st9_b202_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b202_c0 : nS_st8_b202_c1;
  assign nS_st9_b203_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b203_c0 : nS_st8_b203_c1;
  assign nS_st9_b204_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b204_c0 : nS_st8_b204_c1;
  assign nS_st9_b205_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b205_c0 : nS_st8_b205_c1;
  assign nS_st9_b206_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b206_c0 : nS_st8_b206_c1;
  assign nS_st9_b207_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b207_c0 : nS_st8_b207_c1;
  assign nS_st9_b208_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b208_c0 : nS_st8_b208_c1;
  assign nS_st9_b209_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b209_c0 : nS_st8_b209_c1;
  assign nS_st9_b210_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b210_c0 : nS_st8_b210_c1;
  assign nS_st9_b211_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b211_c0 : nS_st8_b211_c1;
  assign nS_st9_b212_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b212_c0 : nS_st8_b212_c1;
  assign nS_st9_b213_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b213_c0 : nS_st8_b213_c1;
  assign nS_st9_b214_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b214_c0 : nS_st8_b214_c1;
  assign nS_st9_b215_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b215_c0 : nS_st8_b215_c1;
  assign nS_st9_b216_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b216_c0 : nS_st8_b216_c1;
  assign nS_st9_b217_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b217_c0 : nS_st8_b217_c1;
  assign nS_st9_b218_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b218_c0 : nS_st8_b218_c1;
  assign nS_st9_b219_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b219_c0 : nS_st8_b219_c1;
  assign nS_st9_b220_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b220_c0 : nS_st8_b220_c1;
  assign nS_st9_b221_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b221_c0 : nS_st8_b221_c1;
  assign nS_st9_b222_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b222_c0 : nS_st8_b222_c1;
  assign nS_st9_b223_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b223_c0 : nS_st8_b223_c1;
  assign nS_st9_b224_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b224_c0 : nS_st8_b224_c1;
  assign nS_st9_b225_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b225_c0 : nS_st8_b225_c1;
  assign nS_st9_b226_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b226_c0 : nS_st8_b226_c1;
  assign nS_st9_b227_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b227_c0 : nS_st8_b227_c1;
  assign nS_st9_b228_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b228_c0 : nS_st8_b228_c1;
  assign nS_st9_b229_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b229_c0 : nS_st8_b229_c1;
  assign nS_st9_b230_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b230_c0 : nS_st8_b230_c1;
  assign nS_st9_b231_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b231_c0 : nS_st8_b231_c1;
  assign nS_st9_b232_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b232_c0 : nS_st8_b232_c1;
  assign nS_st9_b233_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b233_c0 : nS_st8_b233_c1;
  assign nS_st9_b234_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b234_c0 : nS_st8_b234_c1;
  assign nS_st9_b235_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b235_c0 : nS_st8_b235_c1;
  assign nS_st9_b236_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b236_c0 : nS_st8_b236_c1;
  assign nS_st9_b237_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b237_c0 : nS_st8_b237_c1;
  assign nS_st9_b238_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b238_c0 : nS_st8_b238_c1;
  assign nS_st9_b239_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b239_c0 : nS_st8_b239_c1;
  assign nS_st9_b240_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b240_c0 : nS_st8_b240_c1;
  assign nS_st9_b241_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b241_c0 : nS_st8_b241_c1;
  assign nS_st9_b242_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b242_c0 : nS_st8_b242_c1;
  assign nS_st9_b243_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b243_c0 : nS_st8_b243_c1;
  assign nS_st9_b244_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b244_c0 : nS_st8_b244_c1;
  assign nS_st9_b245_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b245_c0 : nS_st8_b245_c1;
  assign nS_st9_b246_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b246_c0 : nS_st8_b246_c1;
  assign nS_st9_b247_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b247_c0 : nS_st8_b247_c1;
  assign nS_st9_b248_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b248_c0 : nS_st8_b248_c1;
  assign nS_st9_b249_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b249_c0 : nS_st8_b249_c1;
  assign nS_st9_b250_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b250_c0 : nS_st8_b250_c1;
  assign nS_st9_b251_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b251_c0 : nS_st8_b251_c1;
  assign nS_st9_b252_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b252_c0 : nS_st8_b252_c1;
  assign nS_st9_b253_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b253_c0 : nS_st8_b253_c1;
  assign nS_st9_b254_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b254_c0 : nS_st8_b254_c1;
  assign nS_st9_b255_c1 = (nC_st8_b127_c1 == 0) ? nS_st8_b255_c0 : nS_st8_b255_c1;
  assign nC_st9_b255_c0 = (nC_st8_b127_c0 == 0) ? nC_st8_b255_c0 : nC_st8_b255_c1;
  assign nC_st9_b255_c1 = (nC_st8_b127_c1 == 0) ? nC_st8_b255_c0 : nC_st8_b255_c1;

  assign out_S[0] = (in_CI == 0) ? nS_st9_b0_c0 : nS_st9_b0_c1;
  assign out_S[1] = (in_CI == 0) ? nS_st9_b1_c0 : nS_st9_b1_c1;
  assign out_S[2] = (in_CI == 0) ? nS_st9_b2_c0 : nS_st9_b2_c1;
  assign out_S[3] = (in_CI == 0) ? nS_st9_b3_c0 : nS_st9_b3_c1;
  assign out_S[4] = (in_CI == 0) ? nS_st9_b4_c0 : nS_st9_b4_c1;
  assign out_S[5] = (in_CI == 0) ? nS_st9_b5_c0 : nS_st9_b5_c1;
  assign out_S[6] = (in_CI == 0) ? nS_st9_b6_c0 : nS_st9_b6_c1;
  assign out_S[7] = (in_CI == 0) ? nS_st9_b7_c0 : nS_st9_b7_c1;
  assign out_S[8] = (in_CI == 0) ? nS_st9_b8_c0 : nS_st9_b8_c1;
  assign out_S[9] = (in_CI == 0) ? nS_st9_b9_c0 : nS_st9_b9_c1;
  assign out_S[10] = (in_CI == 0) ? nS_st9_b10_c0 : nS_st9_b10_c1;
  assign out_S[11] = (in_CI == 0) ? nS_st9_b11_c0 : nS_st9_b11_c1;
  assign out_S[12] = (in_CI == 0) ? nS_st9_b12_c0 : nS_st9_b12_c1;
  assign out_S[13] = (in_CI == 0) ? nS_st9_b13_c0 : nS_st9_b13_c1;
  assign out_S[14] = (in_CI == 0) ? nS_st9_b14_c0 : nS_st9_b14_c1;
  assign out_S[15] = (in_CI == 0) ? nS_st9_b15_c0 : nS_st9_b15_c1;
  assign out_S[16] = (in_CI == 0) ? nS_st9_b16_c0 : nS_st9_b16_c1;
  assign out_S[17] = (in_CI == 0) ? nS_st9_b17_c0 : nS_st9_b17_c1;
  assign out_S[18] = (in_CI == 0) ? nS_st9_b18_c0 : nS_st9_b18_c1;
  assign out_S[19] = (in_CI == 0) ? nS_st9_b19_c0 : nS_st9_b19_c1;
  assign out_S[20] = (in_CI == 0) ? nS_st9_b20_c0 : nS_st9_b20_c1;
  assign out_S[21] = (in_CI == 0) ? nS_st9_b21_c0 : nS_st9_b21_c1;
  assign out_S[22] = (in_CI == 0) ? nS_st9_b22_c0 : nS_st9_b22_c1;
  assign out_S[23] = (in_CI == 0) ? nS_st9_b23_c0 : nS_st9_b23_c1;
  assign out_S[24] = (in_CI == 0) ? nS_st9_b24_c0 : nS_st9_b24_c1;
  assign out_S[25] = (in_CI == 0) ? nS_st9_b25_c0 : nS_st9_b25_c1;
  assign out_S[26] = (in_CI == 0) ? nS_st9_b26_c0 : nS_st9_b26_c1;
  assign out_S[27] = (in_CI == 0) ? nS_st9_b27_c0 : nS_st9_b27_c1;
  assign out_S[28] = (in_CI == 0) ? nS_st9_b28_c0 : nS_st9_b28_c1;
  assign out_S[29] = (in_CI == 0) ? nS_st9_b29_c0 : nS_st9_b29_c1;
  assign out_S[30] = (in_CI == 0) ? nS_st9_b30_c0 : nS_st9_b30_c1;
  assign out_S[31] = (in_CI == 0) ? nS_st9_b31_c0 : nS_st9_b31_c1;
  assign out_S[32] = (in_CI == 0) ? nS_st9_b32_c0 : nS_st9_b32_c1;
  assign out_S[33] = (in_CI == 0) ? nS_st9_b33_c0 : nS_st9_b33_c1;
  assign out_S[34] = (in_CI == 0) ? nS_st9_b34_c0 : nS_st9_b34_c1;
  assign out_S[35] = (in_CI == 0) ? nS_st9_b35_c0 : nS_st9_b35_c1;
  assign out_S[36] = (in_CI == 0) ? nS_st9_b36_c0 : nS_st9_b36_c1;
  assign out_S[37] = (in_CI == 0) ? nS_st9_b37_c0 : nS_st9_b37_c1;
  assign out_S[38] = (in_CI == 0) ? nS_st9_b38_c0 : nS_st9_b38_c1;
  assign out_S[39] = (in_CI == 0) ? nS_st9_b39_c0 : nS_st9_b39_c1;
  assign out_S[40] = (in_CI == 0) ? nS_st9_b40_c0 : nS_st9_b40_c1;
  assign out_S[41] = (in_CI == 0) ? nS_st9_b41_c0 : nS_st9_b41_c1;
  assign out_S[42] = (in_CI == 0) ? nS_st9_b42_c0 : nS_st9_b42_c1;
  assign out_S[43] = (in_CI == 0) ? nS_st9_b43_c0 : nS_st9_b43_c1;
  assign out_S[44] = (in_CI == 0) ? nS_st9_b44_c0 : nS_st9_b44_c1;
  assign out_S[45] = (in_CI == 0) ? nS_st9_b45_c0 : nS_st9_b45_c1;
  assign out_S[46] = (in_CI == 0) ? nS_st9_b46_c0 : nS_st9_b46_c1;
  assign out_S[47] = (in_CI == 0) ? nS_st9_b47_c0 : nS_st9_b47_c1;
  assign out_S[48] = (in_CI == 0) ? nS_st9_b48_c0 : nS_st9_b48_c1;
  assign out_S[49] = (in_CI == 0) ? nS_st9_b49_c0 : nS_st9_b49_c1;
  assign out_S[50] = (in_CI == 0) ? nS_st9_b50_c0 : nS_st9_b50_c1;
  assign out_S[51] = (in_CI == 0) ? nS_st9_b51_c0 : nS_st9_b51_c1;
  assign out_S[52] = (in_CI == 0) ? nS_st9_b52_c0 : nS_st9_b52_c1;
  assign out_S[53] = (in_CI == 0) ? nS_st9_b53_c0 : nS_st9_b53_c1;
  assign out_S[54] = (in_CI == 0) ? nS_st9_b54_c0 : nS_st9_b54_c1;
  assign out_S[55] = (in_CI == 0) ? nS_st9_b55_c0 : nS_st9_b55_c1;
  assign out_S[56] = (in_CI == 0) ? nS_st9_b56_c0 : nS_st9_b56_c1;
  assign out_S[57] = (in_CI == 0) ? nS_st9_b57_c0 : nS_st9_b57_c1;
  assign out_S[58] = (in_CI == 0) ? nS_st9_b58_c0 : nS_st9_b58_c1;
  assign out_S[59] = (in_CI == 0) ? nS_st9_b59_c0 : nS_st9_b59_c1;
  assign out_S[60] = (in_CI == 0) ? nS_st9_b60_c0 : nS_st9_b60_c1;
  assign out_S[61] = (in_CI == 0) ? nS_st9_b61_c0 : nS_st9_b61_c1;
  assign out_S[62] = (in_CI == 0) ? nS_st9_b62_c0 : nS_st9_b62_c1;
  assign out_S[63] = (in_CI == 0) ? nS_st9_b63_c0 : nS_st9_b63_c1;
  assign out_S[64] = (in_CI == 0) ? nS_st9_b64_c0 : nS_st9_b64_c1;
  assign out_S[65] = (in_CI == 0) ? nS_st9_b65_c0 : nS_st9_b65_c1;
  assign out_S[66] = (in_CI == 0) ? nS_st9_b66_c0 : nS_st9_b66_c1;
  assign out_S[67] = (in_CI == 0) ? nS_st9_b67_c0 : nS_st9_b67_c1;
  assign out_S[68] = (in_CI == 0) ? nS_st9_b68_c0 : nS_st9_b68_c1;
  assign out_S[69] = (in_CI == 0) ? nS_st9_b69_c0 : nS_st9_b69_c1;
  assign out_S[70] = (in_CI == 0) ? nS_st9_b70_c0 : nS_st9_b70_c1;
  assign out_S[71] = (in_CI == 0) ? nS_st9_b71_c0 : nS_st9_b71_c1;
  assign out_S[72] = (in_CI == 0) ? nS_st9_b72_c0 : nS_st9_b72_c1;
  assign out_S[73] = (in_CI == 0) ? nS_st9_b73_c0 : nS_st9_b73_c1;
  assign out_S[74] = (in_CI == 0) ? nS_st9_b74_c0 : nS_st9_b74_c1;
  assign out_S[75] = (in_CI == 0) ? nS_st9_b75_c0 : nS_st9_b75_c1;
  assign out_S[76] = (in_CI == 0) ? nS_st9_b76_c0 : nS_st9_b76_c1;
  assign out_S[77] = (in_CI == 0) ? nS_st9_b77_c0 : nS_st9_b77_c1;
  assign out_S[78] = (in_CI == 0) ? nS_st9_b78_c0 : nS_st9_b78_c1;
  assign out_S[79] = (in_CI == 0) ? nS_st9_b79_c0 : nS_st9_b79_c1;
  assign out_S[80] = (in_CI == 0) ? nS_st9_b80_c0 : nS_st9_b80_c1;
  assign out_S[81] = (in_CI == 0) ? nS_st9_b81_c0 : nS_st9_b81_c1;
  assign out_S[82] = (in_CI == 0) ? nS_st9_b82_c0 : nS_st9_b82_c1;
  assign out_S[83] = (in_CI == 0) ? nS_st9_b83_c0 : nS_st9_b83_c1;
  assign out_S[84] = (in_CI == 0) ? nS_st9_b84_c0 : nS_st9_b84_c1;
  assign out_S[85] = (in_CI == 0) ? nS_st9_b85_c0 : nS_st9_b85_c1;
  assign out_S[86] = (in_CI == 0) ? nS_st9_b86_c0 : nS_st9_b86_c1;
  assign out_S[87] = (in_CI == 0) ? nS_st9_b87_c0 : nS_st9_b87_c1;
  assign out_S[88] = (in_CI == 0) ? nS_st9_b88_c0 : nS_st9_b88_c1;
  assign out_S[89] = (in_CI == 0) ? nS_st9_b89_c0 : nS_st9_b89_c1;
  assign out_S[90] = (in_CI == 0) ? nS_st9_b90_c0 : nS_st9_b90_c1;
  assign out_S[91] = (in_CI == 0) ? nS_st9_b91_c0 : nS_st9_b91_c1;
  assign out_S[92] = (in_CI == 0) ? nS_st9_b92_c0 : nS_st9_b92_c1;
  assign out_S[93] = (in_CI == 0) ? nS_st9_b93_c0 : nS_st9_b93_c1;
  assign out_S[94] = (in_CI == 0) ? nS_st9_b94_c0 : nS_st9_b94_c1;
  assign out_S[95] = (in_CI == 0) ? nS_st9_b95_c0 : nS_st9_b95_c1;
  assign out_S[96] = (in_CI == 0) ? nS_st9_b96_c0 : nS_st9_b96_c1;
  assign out_S[97] = (in_CI == 0) ? nS_st9_b97_c0 : nS_st9_b97_c1;
  assign out_S[98] = (in_CI == 0) ? nS_st9_b98_c0 : nS_st9_b98_c1;
  assign out_S[99] = (in_CI == 0) ? nS_st9_b99_c0 : nS_st9_b99_c1;
  assign out_S[100] = (in_CI == 0) ? nS_st9_b100_c0 : nS_st9_b100_c1;
  assign out_S[101] = (in_CI == 0) ? nS_st9_b101_c0 : nS_st9_b101_c1;
  assign out_S[102] = (in_CI == 0) ? nS_st9_b102_c0 : nS_st9_b102_c1;
  assign out_S[103] = (in_CI == 0) ? nS_st9_b103_c0 : nS_st9_b103_c1;
  assign out_S[104] = (in_CI == 0) ? nS_st9_b104_c0 : nS_st9_b104_c1;
  assign out_S[105] = (in_CI == 0) ? nS_st9_b105_c0 : nS_st9_b105_c1;
  assign out_S[106] = (in_CI == 0) ? nS_st9_b106_c0 : nS_st9_b106_c1;
  assign out_S[107] = (in_CI == 0) ? nS_st9_b107_c0 : nS_st9_b107_c1;
  assign out_S[108] = (in_CI == 0) ? nS_st9_b108_c0 : nS_st9_b108_c1;
  assign out_S[109] = (in_CI == 0) ? nS_st9_b109_c0 : nS_st9_b109_c1;
  assign out_S[110] = (in_CI == 0) ? nS_st9_b110_c0 : nS_st9_b110_c1;
  assign out_S[111] = (in_CI == 0) ? nS_st9_b111_c0 : nS_st9_b111_c1;
  assign out_S[112] = (in_CI == 0) ? nS_st9_b112_c0 : nS_st9_b112_c1;
  assign out_S[113] = (in_CI == 0) ? nS_st9_b113_c0 : nS_st9_b113_c1;
  assign out_S[114] = (in_CI == 0) ? nS_st9_b114_c0 : nS_st9_b114_c1;
  assign out_S[115] = (in_CI == 0) ? nS_st9_b115_c0 : nS_st9_b115_c1;
  assign out_S[116] = (in_CI == 0) ? nS_st9_b116_c0 : nS_st9_b116_c1;
  assign out_S[117] = (in_CI == 0) ? nS_st9_b117_c0 : nS_st9_b117_c1;
  assign out_S[118] = (in_CI == 0) ? nS_st9_b118_c0 : nS_st9_b118_c1;
  assign out_S[119] = (in_CI == 0) ? nS_st9_b119_c0 : nS_st9_b119_c1;
  assign out_S[120] = (in_CI == 0) ? nS_st9_b120_c0 : nS_st9_b120_c1;
  assign out_S[121] = (in_CI == 0) ? nS_st9_b121_c0 : nS_st9_b121_c1;
  assign out_S[122] = (in_CI == 0) ? nS_st9_b122_c0 : nS_st9_b122_c1;
  assign out_S[123] = (in_CI == 0) ? nS_st9_b123_c0 : nS_st9_b123_c1;
  assign out_S[124] = (in_CI == 0) ? nS_st9_b124_c0 : nS_st9_b124_c1;
  assign out_S[125] = (in_CI == 0) ? nS_st9_b125_c0 : nS_st9_b125_c1;
  assign out_S[126] = (in_CI == 0) ? nS_st9_b126_c0 : nS_st9_b126_c1;
  assign out_S[127] = (in_CI == 0) ? nS_st9_b127_c0 : nS_st9_b127_c1;
  assign out_S[128] = (in_CI == 0) ? nS_st9_b128_c0 : nS_st9_b128_c1;
  assign out_S[129] = (in_CI == 0) ? nS_st9_b129_c0 : nS_st9_b129_c1;
  assign out_S[130] = (in_CI == 0) ? nS_st9_b130_c0 : nS_st9_b130_c1;
  assign out_S[131] = (in_CI == 0) ? nS_st9_b131_c0 : nS_st9_b131_c1;
  assign out_S[132] = (in_CI == 0) ? nS_st9_b132_c0 : nS_st9_b132_c1;
  assign out_S[133] = (in_CI == 0) ? nS_st9_b133_c0 : nS_st9_b133_c1;
  assign out_S[134] = (in_CI == 0) ? nS_st9_b134_c0 : nS_st9_b134_c1;
  assign out_S[135] = (in_CI == 0) ? nS_st9_b135_c0 : nS_st9_b135_c1;
  assign out_S[136] = (in_CI == 0) ? nS_st9_b136_c0 : nS_st9_b136_c1;
  assign out_S[137] = (in_CI == 0) ? nS_st9_b137_c0 : nS_st9_b137_c1;
  assign out_S[138] = (in_CI == 0) ? nS_st9_b138_c0 : nS_st9_b138_c1;
  assign out_S[139] = (in_CI == 0) ? nS_st9_b139_c0 : nS_st9_b139_c1;
  assign out_S[140] = (in_CI == 0) ? nS_st9_b140_c0 : nS_st9_b140_c1;
  assign out_S[141] = (in_CI == 0) ? nS_st9_b141_c0 : nS_st9_b141_c1;
  assign out_S[142] = (in_CI == 0) ? nS_st9_b142_c0 : nS_st9_b142_c1;
  assign out_S[143] = (in_CI == 0) ? nS_st9_b143_c0 : nS_st9_b143_c1;
  assign out_S[144] = (in_CI == 0) ? nS_st9_b144_c0 : nS_st9_b144_c1;
  assign out_S[145] = (in_CI == 0) ? nS_st9_b145_c0 : nS_st9_b145_c1;
  assign out_S[146] = (in_CI == 0) ? nS_st9_b146_c0 : nS_st9_b146_c1;
  assign out_S[147] = (in_CI == 0) ? nS_st9_b147_c0 : nS_st9_b147_c1;
  assign out_S[148] = (in_CI == 0) ? nS_st9_b148_c0 : nS_st9_b148_c1;
  assign out_S[149] = (in_CI == 0) ? nS_st9_b149_c0 : nS_st9_b149_c1;
  assign out_S[150] = (in_CI == 0) ? nS_st9_b150_c0 : nS_st9_b150_c1;
  assign out_S[151] = (in_CI == 0) ? nS_st9_b151_c0 : nS_st9_b151_c1;
  assign out_S[152] = (in_CI == 0) ? nS_st9_b152_c0 : nS_st9_b152_c1;
  assign out_S[153] = (in_CI == 0) ? nS_st9_b153_c0 : nS_st9_b153_c1;
  assign out_S[154] = (in_CI == 0) ? nS_st9_b154_c0 : nS_st9_b154_c1;
  assign out_S[155] = (in_CI == 0) ? nS_st9_b155_c0 : nS_st9_b155_c1;
  assign out_S[156] = (in_CI == 0) ? nS_st9_b156_c0 : nS_st9_b156_c1;
  assign out_S[157] = (in_CI == 0) ? nS_st9_b157_c0 : nS_st9_b157_c1;
  assign out_S[158] = (in_CI == 0) ? nS_st9_b158_c0 : nS_st9_b158_c1;
  assign out_S[159] = (in_CI == 0) ? nS_st9_b159_c0 : nS_st9_b159_c1;
  assign out_S[160] = (in_CI == 0) ? nS_st9_b160_c0 : nS_st9_b160_c1;
  assign out_S[161] = (in_CI == 0) ? nS_st9_b161_c0 : nS_st9_b161_c1;
  assign out_S[162] = (in_CI == 0) ? nS_st9_b162_c0 : nS_st9_b162_c1;
  assign out_S[163] = (in_CI == 0) ? nS_st9_b163_c0 : nS_st9_b163_c1;
  assign out_S[164] = (in_CI == 0) ? nS_st9_b164_c0 : nS_st9_b164_c1;
  assign out_S[165] = (in_CI == 0) ? nS_st9_b165_c0 : nS_st9_b165_c1;
  assign out_S[166] = (in_CI == 0) ? nS_st9_b166_c0 : nS_st9_b166_c1;
  assign out_S[167] = (in_CI == 0) ? nS_st9_b167_c0 : nS_st9_b167_c1;
  assign out_S[168] = (in_CI == 0) ? nS_st9_b168_c0 : nS_st9_b168_c1;
  assign out_S[169] = (in_CI == 0) ? nS_st9_b169_c0 : nS_st9_b169_c1;
  assign out_S[170] = (in_CI == 0) ? nS_st9_b170_c0 : nS_st9_b170_c1;
  assign out_S[171] = (in_CI == 0) ? nS_st9_b171_c0 : nS_st9_b171_c1;
  assign out_S[172] = (in_CI == 0) ? nS_st9_b172_c0 : nS_st9_b172_c1;
  assign out_S[173] = (in_CI == 0) ? nS_st9_b173_c0 : nS_st9_b173_c1;
  assign out_S[174] = (in_CI == 0) ? nS_st9_b174_c0 : nS_st9_b174_c1;
  assign out_S[175] = (in_CI == 0) ? nS_st9_b175_c0 : nS_st9_b175_c1;
  assign out_S[176] = (in_CI == 0) ? nS_st9_b176_c0 : nS_st9_b176_c1;
  assign out_S[177] = (in_CI == 0) ? nS_st9_b177_c0 : nS_st9_b177_c1;
  assign out_S[178] = (in_CI == 0) ? nS_st9_b178_c0 : nS_st9_b178_c1;
  assign out_S[179] = (in_CI == 0) ? nS_st9_b179_c0 : nS_st9_b179_c1;
  assign out_S[180] = (in_CI == 0) ? nS_st9_b180_c0 : nS_st9_b180_c1;
  assign out_S[181] = (in_CI == 0) ? nS_st9_b181_c0 : nS_st9_b181_c1;
  assign out_S[182] = (in_CI == 0) ? nS_st9_b182_c0 : nS_st9_b182_c1;
  assign out_S[183] = (in_CI == 0) ? nS_st9_b183_c0 : nS_st9_b183_c1;
  assign out_S[184] = (in_CI == 0) ? nS_st9_b184_c0 : nS_st9_b184_c1;
  assign out_S[185] = (in_CI == 0) ? nS_st9_b185_c0 : nS_st9_b185_c1;
  assign out_S[186] = (in_CI == 0) ? nS_st9_b186_c0 : nS_st9_b186_c1;
  assign out_S[187] = (in_CI == 0) ? nS_st9_b187_c0 : nS_st9_b187_c1;
  assign out_S[188] = (in_CI == 0) ? nS_st9_b188_c0 : nS_st9_b188_c1;
  assign out_S[189] = (in_CI == 0) ? nS_st9_b189_c0 : nS_st9_b189_c1;
  assign out_S[190] = (in_CI == 0) ? nS_st9_b190_c0 : nS_st9_b190_c1;
  assign out_S[191] = (in_CI == 0) ? nS_st9_b191_c0 : nS_st9_b191_c1;
  assign out_S[192] = (in_CI == 0) ? nS_st9_b192_c0 : nS_st9_b192_c1;
  assign out_S[193] = (in_CI == 0) ? nS_st9_b193_c0 : nS_st9_b193_c1;
  assign out_S[194] = (in_CI == 0) ? nS_st9_b194_c0 : nS_st9_b194_c1;
  assign out_S[195] = (in_CI == 0) ? nS_st9_b195_c0 : nS_st9_b195_c1;
  assign out_S[196] = (in_CI == 0) ? nS_st9_b196_c0 : nS_st9_b196_c1;
  assign out_S[197] = (in_CI == 0) ? nS_st9_b197_c0 : nS_st9_b197_c1;
  assign out_S[198] = (in_CI == 0) ? nS_st9_b198_c0 : nS_st9_b198_c1;
  assign out_S[199] = (in_CI == 0) ? nS_st9_b199_c0 : nS_st9_b199_c1;
  assign out_S[200] = (in_CI == 0) ? nS_st9_b200_c0 : nS_st9_b200_c1;
  assign out_S[201] = (in_CI == 0) ? nS_st9_b201_c0 : nS_st9_b201_c1;
  assign out_S[202] = (in_CI == 0) ? nS_st9_b202_c0 : nS_st9_b202_c1;
  assign out_S[203] = (in_CI == 0) ? nS_st9_b203_c0 : nS_st9_b203_c1;
  assign out_S[204] = (in_CI == 0) ? nS_st9_b204_c0 : nS_st9_b204_c1;
  assign out_S[205] = (in_CI == 0) ? nS_st9_b205_c0 : nS_st9_b205_c1;
  assign out_S[206] = (in_CI == 0) ? nS_st9_b206_c0 : nS_st9_b206_c1;
  assign out_S[207] = (in_CI == 0) ? nS_st9_b207_c0 : nS_st9_b207_c1;
  assign out_S[208] = (in_CI == 0) ? nS_st9_b208_c0 : nS_st9_b208_c1;
  assign out_S[209] = (in_CI == 0) ? nS_st9_b209_c0 : nS_st9_b209_c1;
  assign out_S[210] = (in_CI == 0) ? nS_st9_b210_c0 : nS_st9_b210_c1;
  assign out_S[211] = (in_CI == 0) ? nS_st9_b211_c0 : nS_st9_b211_c1;
  assign out_S[212] = (in_CI == 0) ? nS_st9_b212_c0 : nS_st9_b212_c1;
  assign out_S[213] = (in_CI == 0) ? nS_st9_b213_c0 : nS_st9_b213_c1;
  assign out_S[214] = (in_CI == 0) ? nS_st9_b214_c0 : nS_st9_b214_c1;
  assign out_S[215] = (in_CI == 0) ? nS_st9_b215_c0 : nS_st9_b215_c1;
  assign out_S[216] = (in_CI == 0) ? nS_st9_b216_c0 : nS_st9_b216_c1;
  assign out_S[217] = (in_CI == 0) ? nS_st9_b217_c0 : nS_st9_b217_c1;
  assign out_S[218] = (in_CI == 0) ? nS_st9_b218_c0 : nS_st9_b218_c1;
  assign out_S[219] = (in_CI == 0) ? nS_st9_b219_c0 : nS_st9_b219_c1;
  assign out_S[220] = (in_CI == 0) ? nS_st9_b220_c0 : nS_st9_b220_c1;
  assign out_S[221] = (in_CI == 0) ? nS_st9_b221_c0 : nS_st9_b221_c1;
  assign out_S[222] = (in_CI == 0) ? nS_st9_b222_c0 : nS_st9_b222_c1;
  assign out_S[223] = (in_CI == 0) ? nS_st9_b223_c0 : nS_st9_b223_c1;
  assign out_S[224] = (in_CI == 0) ? nS_st9_b224_c0 : nS_st9_b224_c1;
  assign out_S[225] = (in_CI == 0) ? nS_st9_b225_c0 : nS_st9_b225_c1;
  assign out_S[226] = (in_CI == 0) ? nS_st9_b226_c0 : nS_st9_b226_c1;
  assign out_S[227] = (in_CI == 0) ? nS_st9_b227_c0 : nS_st9_b227_c1;
  assign out_S[228] = (in_CI == 0) ? nS_st9_b228_c0 : nS_st9_b228_c1;
  assign out_S[229] = (in_CI == 0) ? nS_st9_b229_c0 : nS_st9_b229_c1;
  assign out_S[230] = (in_CI == 0) ? nS_st9_b230_c0 : nS_st9_b230_c1;
  assign out_S[231] = (in_CI == 0) ? nS_st9_b231_c0 : nS_st9_b231_c1;
  assign out_S[232] = (in_CI == 0) ? nS_st9_b232_c0 : nS_st9_b232_c1;
  assign out_S[233] = (in_CI == 0) ? nS_st9_b233_c0 : nS_st9_b233_c1;
  assign out_S[234] = (in_CI == 0) ? nS_st9_b234_c0 : nS_st9_b234_c1;
  assign out_S[235] = (in_CI == 0) ? nS_st9_b235_c0 : nS_st9_b235_c1;
  assign out_S[236] = (in_CI == 0) ? nS_st9_b236_c0 : nS_st9_b236_c1;
  assign out_S[237] = (in_CI == 0) ? nS_st9_b237_c0 : nS_st9_b237_c1;
  assign out_S[238] = (in_CI == 0) ? nS_st9_b238_c0 : nS_st9_b238_c1;
  assign out_S[239] = (in_CI == 0) ? nS_st9_b239_c0 : nS_st9_b239_c1;
  assign out_S[240] = (in_CI == 0) ? nS_st9_b240_c0 : nS_st9_b240_c1;
  assign out_S[241] = (in_CI == 0) ? nS_st9_b241_c0 : nS_st9_b241_c1;
  assign out_S[242] = (in_CI == 0) ? nS_st9_b242_c0 : nS_st9_b242_c1;
  assign out_S[243] = (in_CI == 0) ? nS_st9_b243_c0 : nS_st9_b243_c1;
  assign out_S[244] = (in_CI == 0) ? nS_st9_b244_c0 : nS_st9_b244_c1;
  assign out_S[245] = (in_CI == 0) ? nS_st9_b245_c0 : nS_st9_b245_c1;
  assign out_S[246] = (in_CI == 0) ? nS_st9_b246_c0 : nS_st9_b246_c1;
  assign out_S[247] = (in_CI == 0) ? nS_st9_b247_c0 : nS_st9_b247_c1;
  assign out_S[248] = (in_CI == 0) ? nS_st9_b248_c0 : nS_st9_b248_c1;
  assign out_S[249] = (in_CI == 0) ? nS_st9_b249_c0 : nS_st9_b249_c1;
  assign out_S[250] = (in_CI == 0) ? nS_st9_b250_c0 : nS_st9_b250_c1;
  assign out_S[251] = (in_CI == 0) ? nS_st9_b251_c0 : nS_st9_b251_c1;
  assign out_S[252] = (in_CI == 0) ? nS_st9_b252_c0 : nS_st9_b252_c1;
  assign out_S[253] = (in_CI == 0) ? nS_st9_b253_c0 : nS_st9_b253_c1;
  assign out_S[254] = (in_CI == 0) ? nS_st9_b254_c0 : nS_st9_b254_c1;
  assign out_S[255] = (in_CI == 0) ? nS_st9_b255_c0 : nS_st9_b255_c1;
  assign out_CO = (in_CI == 0) ? nC_st9_b255_c0 : nC_st9_b255_c1;
endmodule

