module VHA (in_A, in_B, out_S, out_CO);
  input in_A, in_B;
  output out_S, out_CO;

  assign out_S = in_A ^ in_B;
  assign out_CO = in_A & in_B;
endmodule

module VFA (in_A, in_B, in_CI, out_S, out_CO);
  input in_A, in_B, in_CI;
  output out_S, out_CO;

  assign out_S = in_A ^ in_B ^ in_CI;
  assign out_CO = (in_A & in_B) | (in_B & in_CI) | (in_CI & in_A);
endmodule



module VCondSumAdder_128 (in_A, in_B, in_CI, out_S, out_CO);
  input [127:0] in_A, in_B;
  input in_CI;
  output [127:0] out_S;
  output out_CO;

  VHA U_st1_b0_c0 (.in_A(in_A[0]), .in_B(in_B[0]), .out_S(nS_st1_b0_c0), .out_CO(nC_st1_b0_c0));
  VFA U_st1_b0_c1 (.in_A(in_A[0]), .in_B(in_B[0]), .in_CI(1'b1), .out_S(nS_st1_b0_c1), .out_CO(nC_st1_b0_c1));
  VHA U_st1_b1_c0 (.in_A(in_A[1]), .in_B(in_B[1]), .out_S(nS_st1_b1_c0), .out_CO(nC_st1_b1_c0));
  VFA U_st1_b1_c1 (.in_A(in_A[1]), .in_B(in_B[1]), .in_CI(1'b1), .out_S(nS_st1_b1_c1), .out_CO(nC_st1_b1_c1));
  VHA U_st1_b2_c0 (.in_A(in_A[2]), .in_B(in_B[2]), .out_S(nS_st1_b2_c0), .out_CO(nC_st1_b2_c0));
  VFA U_st1_b2_c1 (.in_A(in_A[2]), .in_B(in_B[2]), .in_CI(1'b1), .out_S(nS_st1_b2_c1), .out_CO(nC_st1_b2_c1));
  VHA U_st1_b3_c0 (.in_A(in_A[3]), .in_B(in_B[3]), .out_S(nS_st1_b3_c0), .out_CO(nC_st1_b3_c0));
  VFA U_st1_b3_c1 (.in_A(in_A[3]), .in_B(in_B[3]), .in_CI(1'b1), .out_S(nS_st1_b3_c1), .out_CO(nC_st1_b3_c1));
  VHA U_st1_b4_c0 (.in_A(in_A[4]), .in_B(in_B[4]), .out_S(nS_st1_b4_c0), .out_CO(nC_st1_b4_c0));
  VFA U_st1_b4_c1 (.in_A(in_A[4]), .in_B(in_B[4]), .in_CI(1'b1), .out_S(nS_st1_b4_c1), .out_CO(nC_st1_b4_c1));
  VHA U_st1_b5_c0 (.in_A(in_A[5]), .in_B(in_B[5]), .out_S(nS_st1_b5_c0), .out_CO(nC_st1_b5_c0));
  VFA U_st1_b5_c1 (.in_A(in_A[5]), .in_B(in_B[5]), .in_CI(1'b1), .out_S(nS_st1_b5_c1), .out_CO(nC_st1_b5_c1));
  VHA U_st1_b6_c0 (.in_A(in_A[6]), .in_B(in_B[6]), .out_S(nS_st1_b6_c0), .out_CO(nC_st1_b6_c0));
  VFA U_st1_b6_c1 (.in_A(in_A[6]), .in_B(in_B[6]), .in_CI(1'b1), .out_S(nS_st1_b6_c1), .out_CO(nC_st1_b6_c1));
  VHA U_st1_b7_c0 (.in_A(in_A[7]), .in_B(in_B[7]), .out_S(nS_st1_b7_c0), .out_CO(nC_st1_b7_c0));
  VFA U_st1_b7_c1 (.in_A(in_A[7]), .in_B(in_B[7]), .in_CI(1'b1), .out_S(nS_st1_b7_c1), .out_CO(nC_st1_b7_c1));
  VHA U_st1_b8_c0 (.in_A(in_A[8]), .in_B(in_B[8]), .out_S(nS_st1_b8_c0), .out_CO(nC_st1_b8_c0));
  VFA U_st1_b8_c1 (.in_A(in_A[8]), .in_B(in_B[8]), .in_CI(1'b1), .out_S(nS_st1_b8_c1), .out_CO(nC_st1_b8_c1));
  VHA U_st1_b9_c0 (.in_A(in_A[9]), .in_B(in_B[9]), .out_S(nS_st1_b9_c0), .out_CO(nC_st1_b9_c0));
  VFA U_st1_b9_c1 (.in_A(in_A[9]), .in_B(in_B[9]), .in_CI(1'b1), .out_S(nS_st1_b9_c1), .out_CO(nC_st1_b9_c1));
  VHA U_st1_b10_c0 (.in_A(in_A[10]), .in_B(in_B[10]), .out_S(nS_st1_b10_c0), .out_CO(nC_st1_b10_c0));
  VFA U_st1_b10_c1 (.in_A(in_A[10]), .in_B(in_B[10]), .in_CI(1'b1), .out_S(nS_st1_b10_c1), .out_CO(nC_st1_b10_c1));
  VHA U_st1_b11_c0 (.in_A(in_A[11]), .in_B(in_B[11]), .out_S(nS_st1_b11_c0), .out_CO(nC_st1_b11_c0));
  VFA U_st1_b11_c1 (.in_A(in_A[11]), .in_B(in_B[11]), .in_CI(1'b1), .out_S(nS_st1_b11_c1), .out_CO(nC_st1_b11_c1));
  VHA U_st1_b12_c0 (.in_A(in_A[12]), .in_B(in_B[12]), .out_S(nS_st1_b12_c0), .out_CO(nC_st1_b12_c0));
  VFA U_st1_b12_c1 (.in_A(in_A[12]), .in_B(in_B[12]), .in_CI(1'b1), .out_S(nS_st1_b12_c1), .out_CO(nC_st1_b12_c1));
  VHA U_st1_b13_c0 (.in_A(in_A[13]), .in_B(in_B[13]), .out_S(nS_st1_b13_c0), .out_CO(nC_st1_b13_c0));
  VFA U_st1_b13_c1 (.in_A(in_A[13]), .in_B(in_B[13]), .in_CI(1'b1), .out_S(nS_st1_b13_c1), .out_CO(nC_st1_b13_c1));
  VHA U_st1_b14_c0 (.in_A(in_A[14]), .in_B(in_B[14]), .out_S(nS_st1_b14_c0), .out_CO(nC_st1_b14_c0));
  VFA U_st1_b14_c1 (.in_A(in_A[14]), .in_B(in_B[14]), .in_CI(1'b1), .out_S(nS_st1_b14_c1), .out_CO(nC_st1_b14_c1));
  VHA U_st1_b15_c0 (.in_A(in_A[15]), .in_B(in_B[15]), .out_S(nS_st1_b15_c0), .out_CO(nC_st1_b15_c0));
  VFA U_st1_b15_c1 (.in_A(in_A[15]), .in_B(in_B[15]), .in_CI(1'b1), .out_S(nS_st1_b15_c1), .out_CO(nC_st1_b15_c1));
  VHA U_st1_b16_c0 (.in_A(in_A[16]), .in_B(in_B[16]), .out_S(nS_st1_b16_c0), .out_CO(nC_st1_b16_c0));
  VFA U_st1_b16_c1 (.in_A(in_A[16]), .in_B(in_B[16]), .in_CI(1'b1), .out_S(nS_st1_b16_c1), .out_CO(nC_st1_b16_c1));
  VHA U_st1_b17_c0 (.in_A(in_A[17]), .in_B(in_B[17]), .out_S(nS_st1_b17_c0), .out_CO(nC_st1_b17_c0));
  VFA U_st1_b17_c1 (.in_A(in_A[17]), .in_B(in_B[17]), .in_CI(1'b1), .out_S(nS_st1_b17_c1), .out_CO(nC_st1_b17_c1));
  VHA U_st1_b18_c0 (.in_A(in_A[18]), .in_B(in_B[18]), .out_S(nS_st1_b18_c0), .out_CO(nC_st1_b18_c0));
  VFA U_st1_b18_c1 (.in_A(in_A[18]), .in_B(in_B[18]), .in_CI(1'b1), .out_S(nS_st1_b18_c1), .out_CO(nC_st1_b18_c1));
  VHA U_st1_b19_c0 (.in_A(in_A[19]), .in_B(in_B[19]), .out_S(nS_st1_b19_c0), .out_CO(nC_st1_b19_c0));
  VFA U_st1_b19_c1 (.in_A(in_A[19]), .in_B(in_B[19]), .in_CI(1'b1), .out_S(nS_st1_b19_c1), .out_CO(nC_st1_b19_c1));
  VHA U_st1_b20_c0 (.in_A(in_A[20]), .in_B(in_B[20]), .out_S(nS_st1_b20_c0), .out_CO(nC_st1_b20_c0));
  VFA U_st1_b20_c1 (.in_A(in_A[20]), .in_B(in_B[20]), .in_CI(1'b1), .out_S(nS_st1_b20_c1), .out_CO(nC_st1_b20_c1));
  VHA U_st1_b21_c0 (.in_A(in_A[21]), .in_B(in_B[21]), .out_S(nS_st1_b21_c0), .out_CO(nC_st1_b21_c0));
  VFA U_st1_b21_c1 (.in_A(in_A[21]), .in_B(in_B[21]), .in_CI(1'b1), .out_S(nS_st1_b21_c1), .out_CO(nC_st1_b21_c1));
  VHA U_st1_b22_c0 (.in_A(in_A[22]), .in_B(in_B[22]), .out_S(nS_st1_b22_c0), .out_CO(nC_st1_b22_c0));
  VFA U_st1_b22_c1 (.in_A(in_A[22]), .in_B(in_B[22]), .in_CI(1'b1), .out_S(nS_st1_b22_c1), .out_CO(nC_st1_b22_c1));
  VHA U_st1_b23_c0 (.in_A(in_A[23]), .in_B(in_B[23]), .out_S(nS_st1_b23_c0), .out_CO(nC_st1_b23_c0));
  VFA U_st1_b23_c1 (.in_A(in_A[23]), .in_B(in_B[23]), .in_CI(1'b1), .out_S(nS_st1_b23_c1), .out_CO(nC_st1_b23_c1));
  VHA U_st1_b24_c0 (.in_A(in_A[24]), .in_B(in_B[24]), .out_S(nS_st1_b24_c0), .out_CO(nC_st1_b24_c0));
  VFA U_st1_b24_c1 (.in_A(in_A[24]), .in_B(in_B[24]), .in_CI(1'b1), .out_S(nS_st1_b24_c1), .out_CO(nC_st1_b24_c1));
  VHA U_st1_b25_c0 (.in_A(in_A[25]), .in_B(in_B[25]), .out_S(nS_st1_b25_c0), .out_CO(nC_st1_b25_c0));
  VFA U_st1_b25_c1 (.in_A(in_A[25]), .in_B(in_B[25]), .in_CI(1'b1), .out_S(nS_st1_b25_c1), .out_CO(nC_st1_b25_c1));
  VHA U_st1_b26_c0 (.in_A(in_A[26]), .in_B(in_B[26]), .out_S(nS_st1_b26_c0), .out_CO(nC_st1_b26_c0));
  VFA U_st1_b26_c1 (.in_A(in_A[26]), .in_B(in_B[26]), .in_CI(1'b1), .out_S(nS_st1_b26_c1), .out_CO(nC_st1_b26_c1));
  VHA U_st1_b27_c0 (.in_A(in_A[27]), .in_B(in_B[27]), .out_S(nS_st1_b27_c0), .out_CO(nC_st1_b27_c0));
  VFA U_st1_b27_c1 (.in_A(in_A[27]), .in_B(in_B[27]), .in_CI(1'b1), .out_S(nS_st1_b27_c1), .out_CO(nC_st1_b27_c1));
  VHA U_st1_b28_c0 (.in_A(in_A[28]), .in_B(in_B[28]), .out_S(nS_st1_b28_c0), .out_CO(nC_st1_b28_c0));
  VFA U_st1_b28_c1 (.in_A(in_A[28]), .in_B(in_B[28]), .in_CI(1'b1), .out_S(nS_st1_b28_c1), .out_CO(nC_st1_b28_c1));
  VHA U_st1_b29_c0 (.in_A(in_A[29]), .in_B(in_B[29]), .out_S(nS_st1_b29_c0), .out_CO(nC_st1_b29_c0));
  VFA U_st1_b29_c1 (.in_A(in_A[29]), .in_B(in_B[29]), .in_CI(1'b1), .out_S(nS_st1_b29_c1), .out_CO(nC_st1_b29_c1));
  VHA U_st1_b30_c0 (.in_A(in_A[30]), .in_B(in_B[30]), .out_S(nS_st1_b30_c0), .out_CO(nC_st1_b30_c0));
  VFA U_st1_b30_c1 (.in_A(in_A[30]), .in_B(in_B[30]), .in_CI(1'b1), .out_S(nS_st1_b30_c1), .out_CO(nC_st1_b30_c1));
  VHA U_st1_b31_c0 (.in_A(in_A[31]), .in_B(in_B[31]), .out_S(nS_st1_b31_c0), .out_CO(nC_st1_b31_c0));
  VFA U_st1_b31_c1 (.in_A(in_A[31]), .in_B(in_B[31]), .in_CI(1'b1), .out_S(nS_st1_b31_c1), .out_CO(nC_st1_b31_c1));
  VHA U_st1_b32_c0 (.in_A(in_A[32]), .in_B(in_B[32]), .out_S(nS_st1_b32_c0), .out_CO(nC_st1_b32_c0));
  VFA U_st1_b32_c1 (.in_A(in_A[32]), .in_B(in_B[32]), .in_CI(1'b1), .out_S(nS_st1_b32_c1), .out_CO(nC_st1_b32_c1));
  VHA U_st1_b33_c0 (.in_A(in_A[33]), .in_B(in_B[33]), .out_S(nS_st1_b33_c0), .out_CO(nC_st1_b33_c0));
  VFA U_st1_b33_c1 (.in_A(in_A[33]), .in_B(in_B[33]), .in_CI(1'b1), .out_S(nS_st1_b33_c1), .out_CO(nC_st1_b33_c1));
  VHA U_st1_b34_c0 (.in_A(in_A[34]), .in_B(in_B[34]), .out_S(nS_st1_b34_c0), .out_CO(nC_st1_b34_c0));
  VFA U_st1_b34_c1 (.in_A(in_A[34]), .in_B(in_B[34]), .in_CI(1'b1), .out_S(nS_st1_b34_c1), .out_CO(nC_st1_b34_c1));
  VHA U_st1_b35_c0 (.in_A(in_A[35]), .in_B(in_B[35]), .out_S(nS_st1_b35_c0), .out_CO(nC_st1_b35_c0));
  VFA U_st1_b35_c1 (.in_A(in_A[35]), .in_B(in_B[35]), .in_CI(1'b1), .out_S(nS_st1_b35_c1), .out_CO(nC_st1_b35_c1));
  VHA U_st1_b36_c0 (.in_A(in_A[36]), .in_B(in_B[36]), .out_S(nS_st1_b36_c0), .out_CO(nC_st1_b36_c0));
  VFA U_st1_b36_c1 (.in_A(in_A[36]), .in_B(in_B[36]), .in_CI(1'b1), .out_S(nS_st1_b36_c1), .out_CO(nC_st1_b36_c1));
  VHA U_st1_b37_c0 (.in_A(in_A[37]), .in_B(in_B[37]), .out_S(nS_st1_b37_c0), .out_CO(nC_st1_b37_c0));
  VFA U_st1_b37_c1 (.in_A(in_A[37]), .in_B(in_B[37]), .in_CI(1'b1), .out_S(nS_st1_b37_c1), .out_CO(nC_st1_b37_c1));
  VHA U_st1_b38_c0 (.in_A(in_A[38]), .in_B(in_B[38]), .out_S(nS_st1_b38_c0), .out_CO(nC_st1_b38_c0));
  VFA U_st1_b38_c1 (.in_A(in_A[38]), .in_B(in_B[38]), .in_CI(1'b1), .out_S(nS_st1_b38_c1), .out_CO(nC_st1_b38_c1));
  VHA U_st1_b39_c0 (.in_A(in_A[39]), .in_B(in_B[39]), .out_S(nS_st1_b39_c0), .out_CO(nC_st1_b39_c0));
  VFA U_st1_b39_c1 (.in_A(in_A[39]), .in_B(in_B[39]), .in_CI(1'b1), .out_S(nS_st1_b39_c1), .out_CO(nC_st1_b39_c1));
  VHA U_st1_b40_c0 (.in_A(in_A[40]), .in_B(in_B[40]), .out_S(nS_st1_b40_c0), .out_CO(nC_st1_b40_c0));
  VFA U_st1_b40_c1 (.in_A(in_A[40]), .in_B(in_B[40]), .in_CI(1'b1), .out_S(nS_st1_b40_c1), .out_CO(nC_st1_b40_c1));
  VHA U_st1_b41_c0 (.in_A(in_A[41]), .in_B(in_B[41]), .out_S(nS_st1_b41_c0), .out_CO(nC_st1_b41_c0));
  VFA U_st1_b41_c1 (.in_A(in_A[41]), .in_B(in_B[41]), .in_CI(1'b1), .out_S(nS_st1_b41_c1), .out_CO(nC_st1_b41_c1));
  VHA U_st1_b42_c0 (.in_A(in_A[42]), .in_B(in_B[42]), .out_S(nS_st1_b42_c0), .out_CO(nC_st1_b42_c0));
  VFA U_st1_b42_c1 (.in_A(in_A[42]), .in_B(in_B[42]), .in_CI(1'b1), .out_S(nS_st1_b42_c1), .out_CO(nC_st1_b42_c1));
  VHA U_st1_b43_c0 (.in_A(in_A[43]), .in_B(in_B[43]), .out_S(nS_st1_b43_c0), .out_CO(nC_st1_b43_c0));
  VFA U_st1_b43_c1 (.in_A(in_A[43]), .in_B(in_B[43]), .in_CI(1'b1), .out_S(nS_st1_b43_c1), .out_CO(nC_st1_b43_c1));
  VHA U_st1_b44_c0 (.in_A(in_A[44]), .in_B(in_B[44]), .out_S(nS_st1_b44_c0), .out_CO(nC_st1_b44_c0));
  VFA U_st1_b44_c1 (.in_A(in_A[44]), .in_B(in_B[44]), .in_CI(1'b1), .out_S(nS_st1_b44_c1), .out_CO(nC_st1_b44_c1));
  VHA U_st1_b45_c0 (.in_A(in_A[45]), .in_B(in_B[45]), .out_S(nS_st1_b45_c0), .out_CO(nC_st1_b45_c0));
  VFA U_st1_b45_c1 (.in_A(in_A[45]), .in_B(in_B[45]), .in_CI(1'b1), .out_S(nS_st1_b45_c1), .out_CO(nC_st1_b45_c1));
  VHA U_st1_b46_c0 (.in_A(in_A[46]), .in_B(in_B[46]), .out_S(nS_st1_b46_c0), .out_CO(nC_st1_b46_c0));
  VFA U_st1_b46_c1 (.in_A(in_A[46]), .in_B(in_B[46]), .in_CI(1'b1), .out_S(nS_st1_b46_c1), .out_CO(nC_st1_b46_c1));
  VHA U_st1_b47_c0 (.in_A(in_A[47]), .in_B(in_B[47]), .out_S(nS_st1_b47_c0), .out_CO(nC_st1_b47_c0));
  VFA U_st1_b47_c1 (.in_A(in_A[47]), .in_B(in_B[47]), .in_CI(1'b1), .out_S(nS_st1_b47_c1), .out_CO(nC_st1_b47_c1));
  VHA U_st1_b48_c0 (.in_A(in_A[48]), .in_B(in_B[48]), .out_S(nS_st1_b48_c0), .out_CO(nC_st1_b48_c0));
  VFA U_st1_b48_c1 (.in_A(in_A[48]), .in_B(in_B[48]), .in_CI(1'b1), .out_S(nS_st1_b48_c1), .out_CO(nC_st1_b48_c1));
  VHA U_st1_b49_c0 (.in_A(in_A[49]), .in_B(in_B[49]), .out_S(nS_st1_b49_c0), .out_CO(nC_st1_b49_c0));
  VFA U_st1_b49_c1 (.in_A(in_A[49]), .in_B(in_B[49]), .in_CI(1'b1), .out_S(nS_st1_b49_c1), .out_CO(nC_st1_b49_c1));
  VHA U_st1_b50_c0 (.in_A(in_A[50]), .in_B(in_B[50]), .out_S(nS_st1_b50_c0), .out_CO(nC_st1_b50_c0));
  VFA U_st1_b50_c1 (.in_A(in_A[50]), .in_B(in_B[50]), .in_CI(1'b1), .out_S(nS_st1_b50_c1), .out_CO(nC_st1_b50_c1));
  VHA U_st1_b51_c0 (.in_A(in_A[51]), .in_B(in_B[51]), .out_S(nS_st1_b51_c0), .out_CO(nC_st1_b51_c0));
  VFA U_st1_b51_c1 (.in_A(in_A[51]), .in_B(in_B[51]), .in_CI(1'b1), .out_S(nS_st1_b51_c1), .out_CO(nC_st1_b51_c1));
  VHA U_st1_b52_c0 (.in_A(in_A[52]), .in_B(in_B[52]), .out_S(nS_st1_b52_c0), .out_CO(nC_st1_b52_c0));
  VFA U_st1_b52_c1 (.in_A(in_A[52]), .in_B(in_B[52]), .in_CI(1'b1), .out_S(nS_st1_b52_c1), .out_CO(nC_st1_b52_c1));
  VHA U_st1_b53_c0 (.in_A(in_A[53]), .in_B(in_B[53]), .out_S(nS_st1_b53_c0), .out_CO(nC_st1_b53_c0));
  VFA U_st1_b53_c1 (.in_A(in_A[53]), .in_B(in_B[53]), .in_CI(1'b1), .out_S(nS_st1_b53_c1), .out_CO(nC_st1_b53_c1));
  VHA U_st1_b54_c0 (.in_A(in_A[54]), .in_B(in_B[54]), .out_S(nS_st1_b54_c0), .out_CO(nC_st1_b54_c0));
  VFA U_st1_b54_c1 (.in_A(in_A[54]), .in_B(in_B[54]), .in_CI(1'b1), .out_S(nS_st1_b54_c1), .out_CO(nC_st1_b54_c1));
  VHA U_st1_b55_c0 (.in_A(in_A[55]), .in_B(in_B[55]), .out_S(nS_st1_b55_c0), .out_CO(nC_st1_b55_c0));
  VFA U_st1_b55_c1 (.in_A(in_A[55]), .in_B(in_B[55]), .in_CI(1'b1), .out_S(nS_st1_b55_c1), .out_CO(nC_st1_b55_c1));
  VHA U_st1_b56_c0 (.in_A(in_A[56]), .in_B(in_B[56]), .out_S(nS_st1_b56_c0), .out_CO(nC_st1_b56_c0));
  VFA U_st1_b56_c1 (.in_A(in_A[56]), .in_B(in_B[56]), .in_CI(1'b1), .out_S(nS_st1_b56_c1), .out_CO(nC_st1_b56_c1));
  VHA U_st1_b57_c0 (.in_A(in_A[57]), .in_B(in_B[57]), .out_S(nS_st1_b57_c0), .out_CO(nC_st1_b57_c0));
  VFA U_st1_b57_c1 (.in_A(in_A[57]), .in_B(in_B[57]), .in_CI(1'b1), .out_S(nS_st1_b57_c1), .out_CO(nC_st1_b57_c1));
  VHA U_st1_b58_c0 (.in_A(in_A[58]), .in_B(in_B[58]), .out_S(nS_st1_b58_c0), .out_CO(nC_st1_b58_c0));
  VFA U_st1_b58_c1 (.in_A(in_A[58]), .in_B(in_B[58]), .in_CI(1'b1), .out_S(nS_st1_b58_c1), .out_CO(nC_st1_b58_c1));
  VHA U_st1_b59_c0 (.in_A(in_A[59]), .in_B(in_B[59]), .out_S(nS_st1_b59_c0), .out_CO(nC_st1_b59_c0));
  VFA U_st1_b59_c1 (.in_A(in_A[59]), .in_B(in_B[59]), .in_CI(1'b1), .out_S(nS_st1_b59_c1), .out_CO(nC_st1_b59_c1));
  VHA U_st1_b60_c0 (.in_A(in_A[60]), .in_B(in_B[60]), .out_S(nS_st1_b60_c0), .out_CO(nC_st1_b60_c0));
  VFA U_st1_b60_c1 (.in_A(in_A[60]), .in_B(in_B[60]), .in_CI(1'b1), .out_S(nS_st1_b60_c1), .out_CO(nC_st1_b60_c1));
  VHA U_st1_b61_c0 (.in_A(in_A[61]), .in_B(in_B[61]), .out_S(nS_st1_b61_c0), .out_CO(nC_st1_b61_c0));
  VFA U_st1_b61_c1 (.in_A(in_A[61]), .in_B(in_B[61]), .in_CI(1'b1), .out_S(nS_st1_b61_c1), .out_CO(nC_st1_b61_c1));
  VHA U_st1_b62_c0 (.in_A(in_A[62]), .in_B(in_B[62]), .out_S(nS_st1_b62_c0), .out_CO(nC_st1_b62_c0));
  VFA U_st1_b62_c1 (.in_A(in_A[62]), .in_B(in_B[62]), .in_CI(1'b1), .out_S(nS_st1_b62_c1), .out_CO(nC_st1_b62_c1));
  VHA U_st1_b63_c0 (.in_A(in_A[63]), .in_B(in_B[63]), .out_S(nS_st1_b63_c0), .out_CO(nC_st1_b63_c0));
  VFA U_st1_b63_c1 (.in_A(in_A[63]), .in_B(in_B[63]), .in_CI(1'b1), .out_S(nS_st1_b63_c1), .out_CO(nC_st1_b63_c1));
  VHA U_st1_b64_c0 (.in_A(in_A[64]), .in_B(in_B[64]), .out_S(nS_st1_b64_c0), .out_CO(nC_st1_b64_c0));
  VFA U_st1_b64_c1 (.in_A(in_A[64]), .in_B(in_B[64]), .in_CI(1'b1), .out_S(nS_st1_b64_c1), .out_CO(nC_st1_b64_c1));
  VHA U_st1_b65_c0 (.in_A(in_A[65]), .in_B(in_B[65]), .out_S(nS_st1_b65_c0), .out_CO(nC_st1_b65_c0));
  VFA U_st1_b65_c1 (.in_A(in_A[65]), .in_B(in_B[65]), .in_CI(1'b1), .out_S(nS_st1_b65_c1), .out_CO(nC_st1_b65_c1));
  VHA U_st1_b66_c0 (.in_A(in_A[66]), .in_B(in_B[66]), .out_S(nS_st1_b66_c0), .out_CO(nC_st1_b66_c0));
  VFA U_st1_b66_c1 (.in_A(in_A[66]), .in_B(in_B[66]), .in_CI(1'b1), .out_S(nS_st1_b66_c1), .out_CO(nC_st1_b66_c1));
  VHA U_st1_b67_c0 (.in_A(in_A[67]), .in_B(in_B[67]), .out_S(nS_st1_b67_c0), .out_CO(nC_st1_b67_c0));
  VFA U_st1_b67_c1 (.in_A(in_A[67]), .in_B(in_B[67]), .in_CI(1'b1), .out_S(nS_st1_b67_c1), .out_CO(nC_st1_b67_c1));
  VHA U_st1_b68_c0 (.in_A(in_A[68]), .in_B(in_B[68]), .out_S(nS_st1_b68_c0), .out_CO(nC_st1_b68_c0));
  VFA U_st1_b68_c1 (.in_A(in_A[68]), .in_B(in_B[68]), .in_CI(1'b1), .out_S(nS_st1_b68_c1), .out_CO(nC_st1_b68_c1));
  VHA U_st1_b69_c0 (.in_A(in_A[69]), .in_B(in_B[69]), .out_S(nS_st1_b69_c0), .out_CO(nC_st1_b69_c0));
  VFA U_st1_b69_c1 (.in_A(in_A[69]), .in_B(in_B[69]), .in_CI(1'b1), .out_S(nS_st1_b69_c1), .out_CO(nC_st1_b69_c1));
  VHA U_st1_b70_c0 (.in_A(in_A[70]), .in_B(in_B[70]), .out_S(nS_st1_b70_c0), .out_CO(nC_st1_b70_c0));
  VFA U_st1_b70_c1 (.in_A(in_A[70]), .in_B(in_B[70]), .in_CI(1'b1), .out_S(nS_st1_b70_c1), .out_CO(nC_st1_b70_c1));
  VHA U_st1_b71_c0 (.in_A(in_A[71]), .in_B(in_B[71]), .out_S(nS_st1_b71_c0), .out_CO(nC_st1_b71_c0));
  VFA U_st1_b71_c1 (.in_A(in_A[71]), .in_B(in_B[71]), .in_CI(1'b1), .out_S(nS_st1_b71_c1), .out_CO(nC_st1_b71_c1));
  VHA U_st1_b72_c0 (.in_A(in_A[72]), .in_B(in_B[72]), .out_S(nS_st1_b72_c0), .out_CO(nC_st1_b72_c0));
  VFA U_st1_b72_c1 (.in_A(in_A[72]), .in_B(in_B[72]), .in_CI(1'b1), .out_S(nS_st1_b72_c1), .out_CO(nC_st1_b72_c1));
  VHA U_st1_b73_c0 (.in_A(in_A[73]), .in_B(in_B[73]), .out_S(nS_st1_b73_c0), .out_CO(nC_st1_b73_c0));
  VFA U_st1_b73_c1 (.in_A(in_A[73]), .in_B(in_B[73]), .in_CI(1'b1), .out_S(nS_st1_b73_c1), .out_CO(nC_st1_b73_c1));
  VHA U_st1_b74_c0 (.in_A(in_A[74]), .in_B(in_B[74]), .out_S(nS_st1_b74_c0), .out_CO(nC_st1_b74_c0));
  VFA U_st1_b74_c1 (.in_A(in_A[74]), .in_B(in_B[74]), .in_CI(1'b1), .out_S(nS_st1_b74_c1), .out_CO(nC_st1_b74_c1));
  VHA U_st1_b75_c0 (.in_A(in_A[75]), .in_B(in_B[75]), .out_S(nS_st1_b75_c0), .out_CO(nC_st1_b75_c0));
  VFA U_st1_b75_c1 (.in_A(in_A[75]), .in_B(in_B[75]), .in_CI(1'b1), .out_S(nS_st1_b75_c1), .out_CO(nC_st1_b75_c1));
  VHA U_st1_b76_c0 (.in_A(in_A[76]), .in_B(in_B[76]), .out_S(nS_st1_b76_c0), .out_CO(nC_st1_b76_c0));
  VFA U_st1_b76_c1 (.in_A(in_A[76]), .in_B(in_B[76]), .in_CI(1'b1), .out_S(nS_st1_b76_c1), .out_CO(nC_st1_b76_c1));
  VHA U_st1_b77_c0 (.in_A(in_A[77]), .in_B(in_B[77]), .out_S(nS_st1_b77_c0), .out_CO(nC_st1_b77_c0));
  VFA U_st1_b77_c1 (.in_A(in_A[77]), .in_B(in_B[77]), .in_CI(1'b1), .out_S(nS_st1_b77_c1), .out_CO(nC_st1_b77_c1));
  VHA U_st1_b78_c0 (.in_A(in_A[78]), .in_B(in_B[78]), .out_S(nS_st1_b78_c0), .out_CO(nC_st1_b78_c0));
  VFA U_st1_b78_c1 (.in_A(in_A[78]), .in_B(in_B[78]), .in_CI(1'b1), .out_S(nS_st1_b78_c1), .out_CO(nC_st1_b78_c1));
  VHA U_st1_b79_c0 (.in_A(in_A[79]), .in_B(in_B[79]), .out_S(nS_st1_b79_c0), .out_CO(nC_st1_b79_c0));
  VFA U_st1_b79_c1 (.in_A(in_A[79]), .in_B(in_B[79]), .in_CI(1'b1), .out_S(nS_st1_b79_c1), .out_CO(nC_st1_b79_c1));
  VHA U_st1_b80_c0 (.in_A(in_A[80]), .in_B(in_B[80]), .out_S(nS_st1_b80_c0), .out_CO(nC_st1_b80_c0));
  VFA U_st1_b80_c1 (.in_A(in_A[80]), .in_B(in_B[80]), .in_CI(1'b1), .out_S(nS_st1_b80_c1), .out_CO(nC_st1_b80_c1));
  VHA U_st1_b81_c0 (.in_A(in_A[81]), .in_B(in_B[81]), .out_S(nS_st1_b81_c0), .out_CO(nC_st1_b81_c0));
  VFA U_st1_b81_c1 (.in_A(in_A[81]), .in_B(in_B[81]), .in_CI(1'b1), .out_S(nS_st1_b81_c1), .out_CO(nC_st1_b81_c1));
  VHA U_st1_b82_c0 (.in_A(in_A[82]), .in_B(in_B[82]), .out_S(nS_st1_b82_c0), .out_CO(nC_st1_b82_c0));
  VFA U_st1_b82_c1 (.in_A(in_A[82]), .in_B(in_B[82]), .in_CI(1'b1), .out_S(nS_st1_b82_c1), .out_CO(nC_st1_b82_c1));
  VHA U_st1_b83_c0 (.in_A(in_A[83]), .in_B(in_B[83]), .out_S(nS_st1_b83_c0), .out_CO(nC_st1_b83_c0));
  VFA U_st1_b83_c1 (.in_A(in_A[83]), .in_B(in_B[83]), .in_CI(1'b1), .out_S(nS_st1_b83_c1), .out_CO(nC_st1_b83_c1));
  VHA U_st1_b84_c0 (.in_A(in_A[84]), .in_B(in_B[84]), .out_S(nS_st1_b84_c0), .out_CO(nC_st1_b84_c0));
  VFA U_st1_b84_c1 (.in_A(in_A[84]), .in_B(in_B[84]), .in_CI(1'b1), .out_S(nS_st1_b84_c1), .out_CO(nC_st1_b84_c1));
  VHA U_st1_b85_c0 (.in_A(in_A[85]), .in_B(in_B[85]), .out_S(nS_st1_b85_c0), .out_CO(nC_st1_b85_c0));
  VFA U_st1_b85_c1 (.in_A(in_A[85]), .in_B(in_B[85]), .in_CI(1'b1), .out_S(nS_st1_b85_c1), .out_CO(nC_st1_b85_c1));
  VHA U_st1_b86_c0 (.in_A(in_A[86]), .in_B(in_B[86]), .out_S(nS_st1_b86_c0), .out_CO(nC_st1_b86_c0));
  VFA U_st1_b86_c1 (.in_A(in_A[86]), .in_B(in_B[86]), .in_CI(1'b1), .out_S(nS_st1_b86_c1), .out_CO(nC_st1_b86_c1));
  VHA U_st1_b87_c0 (.in_A(in_A[87]), .in_B(in_B[87]), .out_S(nS_st1_b87_c0), .out_CO(nC_st1_b87_c0));
  VFA U_st1_b87_c1 (.in_A(in_A[87]), .in_B(in_B[87]), .in_CI(1'b1), .out_S(nS_st1_b87_c1), .out_CO(nC_st1_b87_c1));
  VHA U_st1_b88_c0 (.in_A(in_A[88]), .in_B(in_B[88]), .out_S(nS_st1_b88_c0), .out_CO(nC_st1_b88_c0));
  VFA U_st1_b88_c1 (.in_A(in_A[88]), .in_B(in_B[88]), .in_CI(1'b1), .out_S(nS_st1_b88_c1), .out_CO(nC_st1_b88_c1));
  VHA U_st1_b89_c0 (.in_A(in_A[89]), .in_B(in_B[89]), .out_S(nS_st1_b89_c0), .out_CO(nC_st1_b89_c0));
  VFA U_st1_b89_c1 (.in_A(in_A[89]), .in_B(in_B[89]), .in_CI(1'b1), .out_S(nS_st1_b89_c1), .out_CO(nC_st1_b89_c1));
  VHA U_st1_b90_c0 (.in_A(in_A[90]), .in_B(in_B[90]), .out_S(nS_st1_b90_c0), .out_CO(nC_st1_b90_c0));
  VFA U_st1_b90_c1 (.in_A(in_A[90]), .in_B(in_B[90]), .in_CI(1'b1), .out_S(nS_st1_b90_c1), .out_CO(nC_st1_b90_c1));
  VHA U_st1_b91_c0 (.in_A(in_A[91]), .in_B(in_B[91]), .out_S(nS_st1_b91_c0), .out_CO(nC_st1_b91_c0));
  VFA U_st1_b91_c1 (.in_A(in_A[91]), .in_B(in_B[91]), .in_CI(1'b1), .out_S(nS_st1_b91_c1), .out_CO(nC_st1_b91_c1));
  VHA U_st1_b92_c0 (.in_A(in_A[92]), .in_B(in_B[92]), .out_S(nS_st1_b92_c0), .out_CO(nC_st1_b92_c0));
  VFA U_st1_b92_c1 (.in_A(in_A[92]), .in_B(in_B[92]), .in_CI(1'b1), .out_S(nS_st1_b92_c1), .out_CO(nC_st1_b92_c1));
  VHA U_st1_b93_c0 (.in_A(in_A[93]), .in_B(in_B[93]), .out_S(nS_st1_b93_c0), .out_CO(nC_st1_b93_c0));
  VFA U_st1_b93_c1 (.in_A(in_A[93]), .in_B(in_B[93]), .in_CI(1'b1), .out_S(nS_st1_b93_c1), .out_CO(nC_st1_b93_c1));
  VHA U_st1_b94_c0 (.in_A(in_A[94]), .in_B(in_B[94]), .out_S(nS_st1_b94_c0), .out_CO(nC_st1_b94_c0));
  VFA U_st1_b94_c1 (.in_A(in_A[94]), .in_B(in_B[94]), .in_CI(1'b1), .out_S(nS_st1_b94_c1), .out_CO(nC_st1_b94_c1));
  VHA U_st1_b95_c0 (.in_A(in_A[95]), .in_B(in_B[95]), .out_S(nS_st1_b95_c0), .out_CO(nC_st1_b95_c0));
  VFA U_st1_b95_c1 (.in_A(in_A[95]), .in_B(in_B[95]), .in_CI(1'b1), .out_S(nS_st1_b95_c1), .out_CO(nC_st1_b95_c1));
  VHA U_st1_b96_c0 (.in_A(in_A[96]), .in_B(in_B[96]), .out_S(nS_st1_b96_c0), .out_CO(nC_st1_b96_c0));
  VFA U_st1_b96_c1 (.in_A(in_A[96]), .in_B(in_B[96]), .in_CI(1'b1), .out_S(nS_st1_b96_c1), .out_CO(nC_st1_b96_c1));
  VHA U_st1_b97_c0 (.in_A(in_A[97]), .in_B(in_B[97]), .out_S(nS_st1_b97_c0), .out_CO(nC_st1_b97_c0));
  VFA U_st1_b97_c1 (.in_A(in_A[97]), .in_B(in_B[97]), .in_CI(1'b1), .out_S(nS_st1_b97_c1), .out_CO(nC_st1_b97_c1));
  VHA U_st1_b98_c0 (.in_A(in_A[98]), .in_B(in_B[98]), .out_S(nS_st1_b98_c0), .out_CO(nC_st1_b98_c0));
  VFA U_st1_b98_c1 (.in_A(in_A[98]), .in_B(in_B[98]), .in_CI(1'b1), .out_S(nS_st1_b98_c1), .out_CO(nC_st1_b98_c1));
  VHA U_st1_b99_c0 (.in_A(in_A[99]), .in_B(in_B[99]), .out_S(nS_st1_b99_c0), .out_CO(nC_st1_b99_c0));
  VFA U_st1_b99_c1 (.in_A(in_A[99]), .in_B(in_B[99]), .in_CI(1'b1), .out_S(nS_st1_b99_c1), .out_CO(nC_st1_b99_c1));
  VHA U_st1_b100_c0 (.in_A(in_A[100]), .in_B(in_B[100]), .out_S(nS_st1_b100_c0), .out_CO(nC_st1_b100_c0));
  VFA U_st1_b100_c1 (.in_A(in_A[100]), .in_B(in_B[100]), .in_CI(1'b1), .out_S(nS_st1_b100_c1), .out_CO(nC_st1_b100_c1));
  VHA U_st1_b101_c0 (.in_A(in_A[101]), .in_B(in_B[101]), .out_S(nS_st1_b101_c0), .out_CO(nC_st1_b101_c0));
  VFA U_st1_b101_c1 (.in_A(in_A[101]), .in_B(in_B[101]), .in_CI(1'b1), .out_S(nS_st1_b101_c1), .out_CO(nC_st1_b101_c1));
  VHA U_st1_b102_c0 (.in_A(in_A[102]), .in_B(in_B[102]), .out_S(nS_st1_b102_c0), .out_CO(nC_st1_b102_c0));
  VFA U_st1_b102_c1 (.in_A(in_A[102]), .in_B(in_B[102]), .in_CI(1'b1), .out_S(nS_st1_b102_c1), .out_CO(nC_st1_b102_c1));
  VHA U_st1_b103_c0 (.in_A(in_A[103]), .in_B(in_B[103]), .out_S(nS_st1_b103_c0), .out_CO(nC_st1_b103_c0));
  VFA U_st1_b103_c1 (.in_A(in_A[103]), .in_B(in_B[103]), .in_CI(1'b1), .out_S(nS_st1_b103_c1), .out_CO(nC_st1_b103_c1));
  VHA U_st1_b104_c0 (.in_A(in_A[104]), .in_B(in_B[104]), .out_S(nS_st1_b104_c0), .out_CO(nC_st1_b104_c0));
  VFA U_st1_b104_c1 (.in_A(in_A[104]), .in_B(in_B[104]), .in_CI(1'b1), .out_S(nS_st1_b104_c1), .out_CO(nC_st1_b104_c1));
  VHA U_st1_b105_c0 (.in_A(in_A[105]), .in_B(in_B[105]), .out_S(nS_st1_b105_c0), .out_CO(nC_st1_b105_c0));
  VFA U_st1_b105_c1 (.in_A(in_A[105]), .in_B(in_B[105]), .in_CI(1'b1), .out_S(nS_st1_b105_c1), .out_CO(nC_st1_b105_c1));
  VHA U_st1_b106_c0 (.in_A(in_A[106]), .in_B(in_B[106]), .out_S(nS_st1_b106_c0), .out_CO(nC_st1_b106_c0));
  VFA U_st1_b106_c1 (.in_A(in_A[106]), .in_B(in_B[106]), .in_CI(1'b1), .out_S(nS_st1_b106_c1), .out_CO(nC_st1_b106_c1));
  VHA U_st1_b107_c0 (.in_A(in_A[107]), .in_B(in_B[107]), .out_S(nS_st1_b107_c0), .out_CO(nC_st1_b107_c0));
  VFA U_st1_b107_c1 (.in_A(in_A[107]), .in_B(in_B[107]), .in_CI(1'b1), .out_S(nS_st1_b107_c1), .out_CO(nC_st1_b107_c1));
  VHA U_st1_b108_c0 (.in_A(in_A[108]), .in_B(in_B[108]), .out_S(nS_st1_b108_c0), .out_CO(nC_st1_b108_c0));
  VFA U_st1_b108_c1 (.in_A(in_A[108]), .in_B(in_B[108]), .in_CI(1'b1), .out_S(nS_st1_b108_c1), .out_CO(nC_st1_b108_c1));
  VHA U_st1_b109_c0 (.in_A(in_A[109]), .in_B(in_B[109]), .out_S(nS_st1_b109_c0), .out_CO(nC_st1_b109_c0));
  VFA U_st1_b109_c1 (.in_A(in_A[109]), .in_B(in_B[109]), .in_CI(1'b1), .out_S(nS_st1_b109_c1), .out_CO(nC_st1_b109_c1));
  VHA U_st1_b110_c0 (.in_A(in_A[110]), .in_B(in_B[110]), .out_S(nS_st1_b110_c0), .out_CO(nC_st1_b110_c0));
  VFA U_st1_b110_c1 (.in_A(in_A[110]), .in_B(in_B[110]), .in_CI(1'b1), .out_S(nS_st1_b110_c1), .out_CO(nC_st1_b110_c1));
  VHA U_st1_b111_c0 (.in_A(in_A[111]), .in_B(in_B[111]), .out_S(nS_st1_b111_c0), .out_CO(nC_st1_b111_c0));
  VFA U_st1_b111_c1 (.in_A(in_A[111]), .in_B(in_B[111]), .in_CI(1'b1), .out_S(nS_st1_b111_c1), .out_CO(nC_st1_b111_c1));
  VHA U_st1_b112_c0 (.in_A(in_A[112]), .in_B(in_B[112]), .out_S(nS_st1_b112_c0), .out_CO(nC_st1_b112_c0));
  VFA U_st1_b112_c1 (.in_A(in_A[112]), .in_B(in_B[112]), .in_CI(1'b1), .out_S(nS_st1_b112_c1), .out_CO(nC_st1_b112_c1));
  VHA U_st1_b113_c0 (.in_A(in_A[113]), .in_B(in_B[113]), .out_S(nS_st1_b113_c0), .out_CO(nC_st1_b113_c0));
  VFA U_st1_b113_c1 (.in_A(in_A[113]), .in_B(in_B[113]), .in_CI(1'b1), .out_S(nS_st1_b113_c1), .out_CO(nC_st1_b113_c1));
  VHA U_st1_b114_c0 (.in_A(in_A[114]), .in_B(in_B[114]), .out_S(nS_st1_b114_c0), .out_CO(nC_st1_b114_c0));
  VFA U_st1_b114_c1 (.in_A(in_A[114]), .in_B(in_B[114]), .in_CI(1'b1), .out_S(nS_st1_b114_c1), .out_CO(nC_st1_b114_c1));
  VHA U_st1_b115_c0 (.in_A(in_A[115]), .in_B(in_B[115]), .out_S(nS_st1_b115_c0), .out_CO(nC_st1_b115_c0));
  VFA U_st1_b115_c1 (.in_A(in_A[115]), .in_B(in_B[115]), .in_CI(1'b1), .out_S(nS_st1_b115_c1), .out_CO(nC_st1_b115_c1));
  VHA U_st1_b116_c0 (.in_A(in_A[116]), .in_B(in_B[116]), .out_S(nS_st1_b116_c0), .out_CO(nC_st1_b116_c0));
  VFA U_st1_b116_c1 (.in_A(in_A[116]), .in_B(in_B[116]), .in_CI(1'b1), .out_S(nS_st1_b116_c1), .out_CO(nC_st1_b116_c1));
  VHA U_st1_b117_c0 (.in_A(in_A[117]), .in_B(in_B[117]), .out_S(nS_st1_b117_c0), .out_CO(nC_st1_b117_c0));
  VFA U_st1_b117_c1 (.in_A(in_A[117]), .in_B(in_B[117]), .in_CI(1'b1), .out_S(nS_st1_b117_c1), .out_CO(nC_st1_b117_c1));
  VHA U_st1_b118_c0 (.in_A(in_A[118]), .in_B(in_B[118]), .out_S(nS_st1_b118_c0), .out_CO(nC_st1_b118_c0));
  VFA U_st1_b118_c1 (.in_A(in_A[118]), .in_B(in_B[118]), .in_CI(1'b1), .out_S(nS_st1_b118_c1), .out_CO(nC_st1_b118_c1));
  VHA U_st1_b119_c0 (.in_A(in_A[119]), .in_B(in_B[119]), .out_S(nS_st1_b119_c0), .out_CO(nC_st1_b119_c0));
  VFA U_st1_b119_c1 (.in_A(in_A[119]), .in_B(in_B[119]), .in_CI(1'b1), .out_S(nS_st1_b119_c1), .out_CO(nC_st1_b119_c1));
  VHA U_st1_b120_c0 (.in_A(in_A[120]), .in_B(in_B[120]), .out_S(nS_st1_b120_c0), .out_CO(nC_st1_b120_c0));
  VFA U_st1_b120_c1 (.in_A(in_A[120]), .in_B(in_B[120]), .in_CI(1'b1), .out_S(nS_st1_b120_c1), .out_CO(nC_st1_b120_c1));
  VHA U_st1_b121_c0 (.in_A(in_A[121]), .in_B(in_B[121]), .out_S(nS_st1_b121_c0), .out_CO(nC_st1_b121_c0));
  VFA U_st1_b121_c1 (.in_A(in_A[121]), .in_B(in_B[121]), .in_CI(1'b1), .out_S(nS_st1_b121_c1), .out_CO(nC_st1_b121_c1));
  VHA U_st1_b122_c0 (.in_A(in_A[122]), .in_B(in_B[122]), .out_S(nS_st1_b122_c0), .out_CO(nC_st1_b122_c0));
  VFA U_st1_b122_c1 (.in_A(in_A[122]), .in_B(in_B[122]), .in_CI(1'b1), .out_S(nS_st1_b122_c1), .out_CO(nC_st1_b122_c1));
  VHA U_st1_b123_c0 (.in_A(in_A[123]), .in_B(in_B[123]), .out_S(nS_st1_b123_c0), .out_CO(nC_st1_b123_c0));
  VFA U_st1_b123_c1 (.in_A(in_A[123]), .in_B(in_B[123]), .in_CI(1'b1), .out_S(nS_st1_b123_c1), .out_CO(nC_st1_b123_c1));
  VHA U_st1_b124_c0 (.in_A(in_A[124]), .in_B(in_B[124]), .out_S(nS_st1_b124_c0), .out_CO(nC_st1_b124_c0));
  VFA U_st1_b124_c1 (.in_A(in_A[124]), .in_B(in_B[124]), .in_CI(1'b1), .out_S(nS_st1_b124_c1), .out_CO(nC_st1_b124_c1));
  VHA U_st1_b125_c0 (.in_A(in_A[125]), .in_B(in_B[125]), .out_S(nS_st1_b125_c0), .out_CO(nC_st1_b125_c0));
  VFA U_st1_b125_c1 (.in_A(in_A[125]), .in_B(in_B[125]), .in_CI(1'b1), .out_S(nS_st1_b125_c1), .out_CO(nC_st1_b125_c1));
  VHA U_st1_b126_c0 (.in_A(in_A[126]), .in_B(in_B[126]), .out_S(nS_st1_b126_c0), .out_CO(nC_st1_b126_c0));
  VFA U_st1_b126_c1 (.in_A(in_A[126]), .in_B(in_B[126]), .in_CI(1'b1), .out_S(nS_st1_b126_c1), .out_CO(nC_st1_b126_c1));
  VHA U_st1_b127_c0 (.in_A(in_A[127]), .in_B(in_B[127]), .out_S(nS_st1_b127_c0), .out_CO(nC_st1_b127_c0));
  VFA U_st1_b127_c1 (.in_A(in_A[127]), .in_B(in_B[127]), .in_CI(1'b1), .out_S(nS_st1_b127_c1), .out_CO(nC_st1_b127_c1));

  assign nS_st2_b0_c0 = nS_st1_b0_c0;
  assign nS_st2_b1_c0 = (nC_st1_b0_c0 == 0) ? nS_st1_b1_c0 : nS_st1_b1_c1;
  assign nS_st2_b2_c0 = nS_st1_b2_c0;
  assign nS_st2_b3_c0 = (nC_st1_b2_c0 == 0) ? nS_st1_b3_c0 : nS_st1_b3_c1;
  assign nS_st2_b4_c0 = nS_st1_b4_c0;
  assign nS_st2_b5_c0 = (nC_st1_b4_c0 == 0) ? nS_st1_b5_c0 : nS_st1_b5_c1;
  assign nS_st2_b6_c0 = nS_st1_b6_c0;
  assign nS_st2_b7_c0 = (nC_st1_b6_c0 == 0) ? nS_st1_b7_c0 : nS_st1_b7_c1;
  assign nS_st2_b8_c0 = nS_st1_b8_c0;
  assign nS_st2_b9_c0 = (nC_st1_b8_c0 == 0) ? nS_st1_b9_c0 : nS_st1_b9_c1;
  assign nS_st2_b10_c0 = nS_st1_b10_c0;
  assign nS_st2_b11_c0 = (nC_st1_b10_c0 == 0) ? nS_st1_b11_c0 : nS_st1_b11_c1;
  assign nS_st2_b12_c0 = nS_st1_b12_c0;
  assign nS_st2_b13_c0 = (nC_st1_b12_c0 == 0) ? nS_st1_b13_c0 : nS_st1_b13_c1;
  assign nS_st2_b14_c0 = nS_st1_b14_c0;
  assign nS_st2_b15_c0 = (nC_st1_b14_c0 == 0) ? nS_st1_b15_c0 : nS_st1_b15_c1;
  assign nS_st2_b16_c0 = nS_st1_b16_c0;
  assign nS_st2_b17_c0 = (nC_st1_b16_c0 == 0) ? nS_st1_b17_c0 : nS_st1_b17_c1;
  assign nS_st2_b18_c0 = nS_st1_b18_c0;
  assign nS_st2_b19_c0 = (nC_st1_b18_c0 == 0) ? nS_st1_b19_c0 : nS_st1_b19_c1;
  assign nS_st2_b20_c0 = nS_st1_b20_c0;
  assign nS_st2_b21_c0 = (nC_st1_b20_c0 == 0) ? nS_st1_b21_c0 : nS_st1_b21_c1;
  assign nS_st2_b22_c0 = nS_st1_b22_c0;
  assign nS_st2_b23_c0 = (nC_st1_b22_c0 == 0) ? nS_st1_b23_c0 : nS_st1_b23_c1;
  assign nS_st2_b24_c0 = nS_st1_b24_c0;
  assign nS_st2_b25_c0 = (nC_st1_b24_c0 == 0) ? nS_st1_b25_c0 : nS_st1_b25_c1;
  assign nS_st2_b26_c0 = nS_st1_b26_c0;
  assign nS_st2_b27_c0 = (nC_st1_b26_c0 == 0) ? nS_st1_b27_c0 : nS_st1_b27_c1;
  assign nS_st2_b28_c0 = nS_st1_b28_c0;
  assign nS_st2_b29_c0 = (nC_st1_b28_c0 == 0) ? nS_st1_b29_c0 : nS_st1_b29_c1;
  assign nS_st2_b30_c0 = nS_st1_b30_c0;
  assign nS_st2_b31_c0 = (nC_st1_b30_c0 == 0) ? nS_st1_b31_c0 : nS_st1_b31_c1;
  assign nS_st2_b32_c0 = nS_st1_b32_c0;
  assign nS_st2_b33_c0 = (nC_st1_b32_c0 == 0) ? nS_st1_b33_c0 : nS_st1_b33_c1;
  assign nS_st2_b34_c0 = nS_st1_b34_c0;
  assign nS_st2_b35_c0 = (nC_st1_b34_c0 == 0) ? nS_st1_b35_c0 : nS_st1_b35_c1;
  assign nS_st2_b36_c0 = nS_st1_b36_c0;
  assign nS_st2_b37_c0 = (nC_st1_b36_c0 == 0) ? nS_st1_b37_c0 : nS_st1_b37_c1;
  assign nS_st2_b38_c0 = nS_st1_b38_c0;
  assign nS_st2_b39_c0 = (nC_st1_b38_c0 == 0) ? nS_st1_b39_c0 : nS_st1_b39_c1;
  assign nS_st2_b40_c0 = nS_st1_b40_c0;
  assign nS_st2_b41_c0 = (nC_st1_b40_c0 == 0) ? nS_st1_b41_c0 : nS_st1_b41_c1;
  assign nS_st2_b42_c0 = nS_st1_b42_c0;
  assign nS_st2_b43_c0 = (nC_st1_b42_c0 == 0) ? nS_st1_b43_c0 : nS_st1_b43_c1;
  assign nS_st2_b44_c0 = nS_st1_b44_c0;
  assign nS_st2_b45_c0 = (nC_st1_b44_c0 == 0) ? nS_st1_b45_c0 : nS_st1_b45_c1;
  assign nS_st2_b46_c0 = nS_st1_b46_c0;
  assign nS_st2_b47_c0 = (nC_st1_b46_c0 == 0) ? nS_st1_b47_c0 : nS_st1_b47_c1;
  assign nS_st2_b48_c0 = nS_st1_b48_c0;
  assign nS_st2_b49_c0 = (nC_st1_b48_c0 == 0) ? nS_st1_b49_c0 : nS_st1_b49_c1;
  assign nS_st2_b50_c0 = nS_st1_b50_c0;
  assign nS_st2_b51_c0 = (nC_st1_b50_c0 == 0) ? nS_st1_b51_c0 : nS_st1_b51_c1;
  assign nS_st2_b52_c0 = nS_st1_b52_c0;
  assign nS_st2_b53_c0 = (nC_st1_b52_c0 == 0) ? nS_st1_b53_c0 : nS_st1_b53_c1;
  assign nS_st2_b54_c0 = nS_st1_b54_c0;
  assign nS_st2_b55_c0 = (nC_st1_b54_c0 == 0) ? nS_st1_b55_c0 : nS_st1_b55_c1;
  assign nS_st2_b56_c0 = nS_st1_b56_c0;
  assign nS_st2_b57_c0 = (nC_st1_b56_c0 == 0) ? nS_st1_b57_c0 : nS_st1_b57_c1;
  assign nS_st2_b58_c0 = nS_st1_b58_c0;
  assign nS_st2_b59_c0 = (nC_st1_b58_c0 == 0) ? nS_st1_b59_c0 : nS_st1_b59_c1;
  assign nS_st2_b60_c0 = nS_st1_b60_c0;
  assign nS_st2_b61_c0 = (nC_st1_b60_c0 == 0) ? nS_st1_b61_c0 : nS_st1_b61_c1;
  assign nS_st2_b62_c0 = nS_st1_b62_c0;
  assign nS_st2_b63_c0 = (nC_st1_b62_c0 == 0) ? nS_st1_b63_c0 : nS_st1_b63_c1;
  assign nS_st2_b64_c0 = nS_st1_b64_c0;
  assign nS_st2_b65_c0 = (nC_st1_b64_c0 == 0) ? nS_st1_b65_c0 : nS_st1_b65_c1;
  assign nS_st2_b66_c0 = nS_st1_b66_c0;
  assign nS_st2_b67_c0 = (nC_st1_b66_c0 == 0) ? nS_st1_b67_c0 : nS_st1_b67_c1;
  assign nS_st2_b68_c0 = nS_st1_b68_c0;
  assign nS_st2_b69_c0 = (nC_st1_b68_c0 == 0) ? nS_st1_b69_c0 : nS_st1_b69_c1;
  assign nS_st2_b70_c0 = nS_st1_b70_c0;
  assign nS_st2_b71_c0 = (nC_st1_b70_c0 == 0) ? nS_st1_b71_c0 : nS_st1_b71_c1;
  assign nS_st2_b72_c0 = nS_st1_b72_c0;
  assign nS_st2_b73_c0 = (nC_st1_b72_c0 == 0) ? nS_st1_b73_c0 : nS_st1_b73_c1;
  assign nS_st2_b74_c0 = nS_st1_b74_c0;
  assign nS_st2_b75_c0 = (nC_st1_b74_c0 == 0) ? nS_st1_b75_c0 : nS_st1_b75_c1;
  assign nS_st2_b76_c0 = nS_st1_b76_c0;
  assign nS_st2_b77_c0 = (nC_st1_b76_c0 == 0) ? nS_st1_b77_c0 : nS_st1_b77_c1;
  assign nS_st2_b78_c0 = nS_st1_b78_c0;
  assign nS_st2_b79_c0 = (nC_st1_b78_c0 == 0) ? nS_st1_b79_c0 : nS_st1_b79_c1;
  assign nS_st2_b80_c0 = nS_st1_b80_c0;
  assign nS_st2_b81_c0 = (nC_st1_b80_c0 == 0) ? nS_st1_b81_c0 : nS_st1_b81_c1;
  assign nS_st2_b82_c0 = nS_st1_b82_c0;
  assign nS_st2_b83_c0 = (nC_st1_b82_c0 == 0) ? nS_st1_b83_c0 : nS_st1_b83_c1;
  assign nS_st2_b84_c0 = nS_st1_b84_c0;
  assign nS_st2_b85_c0 = (nC_st1_b84_c0 == 0) ? nS_st1_b85_c0 : nS_st1_b85_c1;
  assign nS_st2_b86_c0 = nS_st1_b86_c0;
  assign nS_st2_b87_c0 = (nC_st1_b86_c0 == 0) ? nS_st1_b87_c0 : nS_st1_b87_c1;
  assign nS_st2_b88_c0 = nS_st1_b88_c0;
  assign nS_st2_b89_c0 = (nC_st1_b88_c0 == 0) ? nS_st1_b89_c0 : nS_st1_b89_c1;
  assign nS_st2_b90_c0 = nS_st1_b90_c0;
  assign nS_st2_b91_c0 = (nC_st1_b90_c0 == 0) ? nS_st1_b91_c0 : nS_st1_b91_c1;
  assign nS_st2_b92_c0 = nS_st1_b92_c0;
  assign nS_st2_b93_c0 = (nC_st1_b92_c0 == 0) ? nS_st1_b93_c0 : nS_st1_b93_c1;
  assign nS_st2_b94_c0 = nS_st1_b94_c0;
  assign nS_st2_b95_c0 = (nC_st1_b94_c0 == 0) ? nS_st1_b95_c0 : nS_st1_b95_c1;
  assign nS_st2_b96_c0 = nS_st1_b96_c0;
  assign nS_st2_b97_c0 = (nC_st1_b96_c0 == 0) ? nS_st1_b97_c0 : nS_st1_b97_c1;
  assign nS_st2_b98_c0 = nS_st1_b98_c0;
  assign nS_st2_b99_c0 = (nC_st1_b98_c0 == 0) ? nS_st1_b99_c0 : nS_st1_b99_c1;
  assign nS_st2_b100_c0 = nS_st1_b100_c0;
  assign nS_st2_b101_c0 = (nC_st1_b100_c0 == 0) ? nS_st1_b101_c0 : nS_st1_b101_c1;
  assign nS_st2_b102_c0 = nS_st1_b102_c0;
  assign nS_st2_b103_c0 = (nC_st1_b102_c0 == 0) ? nS_st1_b103_c0 : nS_st1_b103_c1;
  assign nS_st2_b104_c0 = nS_st1_b104_c0;
  assign nS_st2_b105_c0 = (nC_st1_b104_c0 == 0) ? nS_st1_b105_c0 : nS_st1_b105_c1;
  assign nS_st2_b106_c0 = nS_st1_b106_c0;
  assign nS_st2_b107_c0 = (nC_st1_b106_c0 == 0) ? nS_st1_b107_c0 : nS_st1_b107_c1;
  assign nS_st2_b108_c0 = nS_st1_b108_c0;
  assign nS_st2_b109_c0 = (nC_st1_b108_c0 == 0) ? nS_st1_b109_c0 : nS_st1_b109_c1;
  assign nS_st2_b110_c0 = nS_st1_b110_c0;
  assign nS_st2_b111_c0 = (nC_st1_b110_c0 == 0) ? nS_st1_b111_c0 : nS_st1_b111_c1;
  assign nS_st2_b112_c0 = nS_st1_b112_c0;
  assign nS_st2_b113_c0 = (nC_st1_b112_c0 == 0) ? nS_st1_b113_c0 : nS_st1_b113_c1;
  assign nS_st2_b114_c0 = nS_st1_b114_c0;
  assign nS_st2_b115_c0 = (nC_st1_b114_c0 == 0) ? nS_st1_b115_c0 : nS_st1_b115_c1;
  assign nS_st2_b116_c0 = nS_st1_b116_c0;
  assign nS_st2_b117_c0 = (nC_st1_b116_c0 == 0) ? nS_st1_b117_c0 : nS_st1_b117_c1;
  assign nS_st2_b118_c0 = nS_st1_b118_c0;
  assign nS_st2_b119_c0 = (nC_st1_b118_c0 == 0) ? nS_st1_b119_c0 : nS_st1_b119_c1;
  assign nS_st2_b120_c0 = nS_st1_b120_c0;
  assign nS_st2_b121_c0 = (nC_st1_b120_c0 == 0) ? nS_st1_b121_c0 : nS_st1_b121_c1;
  assign nS_st2_b122_c0 = nS_st1_b122_c0;
  assign nS_st2_b123_c0 = (nC_st1_b122_c0 == 0) ? nS_st1_b123_c0 : nS_st1_b123_c1;
  assign nS_st2_b124_c0 = nS_st1_b124_c0;
  assign nS_st2_b125_c0 = (nC_st1_b124_c0 == 0) ? nS_st1_b125_c0 : nS_st1_b125_c1;
  assign nS_st2_b126_c0 = nS_st1_b126_c0;
  assign nS_st2_b127_c0 = (nC_st1_b126_c0 == 0) ? nS_st1_b127_c0 : nS_st1_b127_c1;
  assign nS_st2_b0_c1 = nS_st1_b0_c1;
  assign nS_st2_b1_c1 = (nC_st1_b0_c1 == 0) ? nS_st1_b1_c0 : nS_st1_b1_c1;
  assign nS_st2_b2_c1 = nS_st1_b2_c1;
  assign nS_st2_b3_c1 = (nC_st1_b2_c1 == 0) ? nS_st1_b3_c0 : nS_st1_b3_c1;
  assign nS_st2_b4_c1 = nS_st1_b4_c1;
  assign nS_st2_b5_c1 = (nC_st1_b4_c1 == 0) ? nS_st1_b5_c0 : nS_st1_b5_c1;
  assign nS_st2_b6_c1 = nS_st1_b6_c1;
  assign nS_st2_b7_c1 = (nC_st1_b6_c1 == 0) ? nS_st1_b7_c0 : nS_st1_b7_c1;
  assign nS_st2_b8_c1 = nS_st1_b8_c1;
  assign nS_st2_b9_c1 = (nC_st1_b8_c1 == 0) ? nS_st1_b9_c0 : nS_st1_b9_c1;
  assign nS_st2_b10_c1 = nS_st1_b10_c1;
  assign nS_st2_b11_c1 = (nC_st1_b10_c1 == 0) ? nS_st1_b11_c0 : nS_st1_b11_c1;
  assign nS_st2_b12_c1 = nS_st1_b12_c1;
  assign nS_st2_b13_c1 = (nC_st1_b12_c1 == 0) ? nS_st1_b13_c0 : nS_st1_b13_c1;
  assign nS_st2_b14_c1 = nS_st1_b14_c1;
  assign nS_st2_b15_c1 = (nC_st1_b14_c1 == 0) ? nS_st1_b15_c0 : nS_st1_b15_c1;
  assign nS_st2_b16_c1 = nS_st1_b16_c1;
  assign nS_st2_b17_c1 = (nC_st1_b16_c1 == 0) ? nS_st1_b17_c0 : nS_st1_b17_c1;
  assign nS_st2_b18_c1 = nS_st1_b18_c1;
  assign nS_st2_b19_c1 = (nC_st1_b18_c1 == 0) ? nS_st1_b19_c0 : nS_st1_b19_c1;
  assign nS_st2_b20_c1 = nS_st1_b20_c1;
  assign nS_st2_b21_c1 = (nC_st1_b20_c1 == 0) ? nS_st1_b21_c0 : nS_st1_b21_c1;
  assign nS_st2_b22_c1 = nS_st1_b22_c1;
  assign nS_st2_b23_c1 = (nC_st1_b22_c1 == 0) ? nS_st1_b23_c0 : nS_st1_b23_c1;
  assign nS_st2_b24_c1 = nS_st1_b24_c1;
  assign nS_st2_b25_c1 = (nC_st1_b24_c1 == 0) ? nS_st1_b25_c0 : nS_st1_b25_c1;
  assign nS_st2_b26_c1 = nS_st1_b26_c1;
  assign nS_st2_b27_c1 = (nC_st1_b26_c1 == 0) ? nS_st1_b27_c0 : nS_st1_b27_c1;
  assign nS_st2_b28_c1 = nS_st1_b28_c1;
  assign nS_st2_b29_c1 = (nC_st1_b28_c1 == 0) ? nS_st1_b29_c0 : nS_st1_b29_c1;
  assign nS_st2_b30_c1 = nS_st1_b30_c1;
  assign nS_st2_b31_c1 = (nC_st1_b30_c1 == 0) ? nS_st1_b31_c0 : nS_st1_b31_c1;
  assign nS_st2_b32_c1 = nS_st1_b32_c1;
  assign nS_st2_b33_c1 = (nC_st1_b32_c1 == 0) ? nS_st1_b33_c0 : nS_st1_b33_c1;
  assign nS_st2_b34_c1 = nS_st1_b34_c1;
  assign nS_st2_b35_c1 = (nC_st1_b34_c1 == 0) ? nS_st1_b35_c0 : nS_st1_b35_c1;
  assign nS_st2_b36_c1 = nS_st1_b36_c1;
  assign nS_st2_b37_c1 = (nC_st1_b36_c1 == 0) ? nS_st1_b37_c0 : nS_st1_b37_c1;
  assign nS_st2_b38_c1 = nS_st1_b38_c1;
  assign nS_st2_b39_c1 = (nC_st1_b38_c1 == 0) ? nS_st1_b39_c0 : nS_st1_b39_c1;
  assign nS_st2_b40_c1 = nS_st1_b40_c1;
  assign nS_st2_b41_c1 = (nC_st1_b40_c1 == 0) ? nS_st1_b41_c0 : nS_st1_b41_c1;
  assign nS_st2_b42_c1 = nS_st1_b42_c1;
  assign nS_st2_b43_c1 = (nC_st1_b42_c1 == 0) ? nS_st1_b43_c0 : nS_st1_b43_c1;
  assign nS_st2_b44_c1 = nS_st1_b44_c1;
  assign nS_st2_b45_c1 = (nC_st1_b44_c1 == 0) ? nS_st1_b45_c0 : nS_st1_b45_c1;
  assign nS_st2_b46_c1 = nS_st1_b46_c1;
  assign nS_st2_b47_c1 = (nC_st1_b46_c1 == 0) ? nS_st1_b47_c0 : nS_st1_b47_c1;
  assign nS_st2_b48_c1 = nS_st1_b48_c1;
  assign nS_st2_b49_c1 = (nC_st1_b48_c1 == 0) ? nS_st1_b49_c0 : nS_st1_b49_c1;
  assign nS_st2_b50_c1 = nS_st1_b50_c1;
  assign nS_st2_b51_c1 = (nC_st1_b50_c1 == 0) ? nS_st1_b51_c0 : nS_st1_b51_c1;
  assign nS_st2_b52_c1 = nS_st1_b52_c1;
  assign nS_st2_b53_c1 = (nC_st1_b52_c1 == 0) ? nS_st1_b53_c0 : nS_st1_b53_c1;
  assign nS_st2_b54_c1 = nS_st1_b54_c1;
  assign nS_st2_b55_c1 = (nC_st1_b54_c1 == 0) ? nS_st1_b55_c0 : nS_st1_b55_c1;
  assign nS_st2_b56_c1 = nS_st1_b56_c1;
  assign nS_st2_b57_c1 = (nC_st1_b56_c1 == 0) ? nS_st1_b57_c0 : nS_st1_b57_c1;
  assign nS_st2_b58_c1 = nS_st1_b58_c1;
  assign nS_st2_b59_c1 = (nC_st1_b58_c1 == 0) ? nS_st1_b59_c0 : nS_st1_b59_c1;
  assign nS_st2_b60_c1 = nS_st1_b60_c1;
  assign nS_st2_b61_c1 = (nC_st1_b60_c1 == 0) ? nS_st1_b61_c0 : nS_st1_b61_c1;
  assign nS_st2_b62_c1 = nS_st1_b62_c1;
  assign nS_st2_b63_c1 = (nC_st1_b62_c1 == 0) ? nS_st1_b63_c0 : nS_st1_b63_c1;
  assign nS_st2_b64_c1 = nS_st1_b64_c1;
  assign nS_st2_b65_c1 = (nC_st1_b64_c1 == 0) ? nS_st1_b65_c0 : nS_st1_b65_c1;
  assign nS_st2_b66_c1 = nS_st1_b66_c1;
  assign nS_st2_b67_c1 = (nC_st1_b66_c1 == 0) ? nS_st1_b67_c0 : nS_st1_b67_c1;
  assign nS_st2_b68_c1 = nS_st1_b68_c1;
  assign nS_st2_b69_c1 = (nC_st1_b68_c1 == 0) ? nS_st1_b69_c0 : nS_st1_b69_c1;
  assign nS_st2_b70_c1 = nS_st1_b70_c1;
  assign nS_st2_b71_c1 = (nC_st1_b70_c1 == 0) ? nS_st1_b71_c0 : nS_st1_b71_c1;
  assign nS_st2_b72_c1 = nS_st1_b72_c1;
  assign nS_st2_b73_c1 = (nC_st1_b72_c1 == 0) ? nS_st1_b73_c0 : nS_st1_b73_c1;
  assign nS_st2_b74_c1 = nS_st1_b74_c1;
  assign nS_st2_b75_c1 = (nC_st1_b74_c1 == 0) ? nS_st1_b75_c0 : nS_st1_b75_c1;
  assign nS_st2_b76_c1 = nS_st1_b76_c1;
  assign nS_st2_b77_c1 = (nC_st1_b76_c1 == 0) ? nS_st1_b77_c0 : nS_st1_b77_c1;
  assign nS_st2_b78_c1 = nS_st1_b78_c1;
  assign nS_st2_b79_c1 = (nC_st1_b78_c1 == 0) ? nS_st1_b79_c0 : nS_st1_b79_c1;
  assign nS_st2_b80_c1 = nS_st1_b80_c1;
  assign nS_st2_b81_c1 = (nC_st1_b80_c1 == 0) ? nS_st1_b81_c0 : nS_st1_b81_c1;
  assign nS_st2_b82_c1 = nS_st1_b82_c1;
  assign nS_st2_b83_c1 = (nC_st1_b82_c1 == 0) ? nS_st1_b83_c0 : nS_st1_b83_c1;
  assign nS_st2_b84_c1 = nS_st1_b84_c1;
  assign nS_st2_b85_c1 = (nC_st1_b84_c1 == 0) ? nS_st1_b85_c0 : nS_st1_b85_c1;
  assign nS_st2_b86_c1 = nS_st1_b86_c1;
  assign nS_st2_b87_c1 = (nC_st1_b86_c1 == 0) ? nS_st1_b87_c0 : nS_st1_b87_c1;
  assign nS_st2_b88_c1 = nS_st1_b88_c1;
  assign nS_st2_b89_c1 = (nC_st1_b88_c1 == 0) ? nS_st1_b89_c0 : nS_st1_b89_c1;
  assign nS_st2_b90_c1 = nS_st1_b90_c1;
  assign nS_st2_b91_c1 = (nC_st1_b90_c1 == 0) ? nS_st1_b91_c0 : nS_st1_b91_c1;
  assign nS_st2_b92_c1 = nS_st1_b92_c1;
  assign nS_st2_b93_c1 = (nC_st1_b92_c1 == 0) ? nS_st1_b93_c0 : nS_st1_b93_c1;
  assign nS_st2_b94_c1 = nS_st1_b94_c1;
  assign nS_st2_b95_c1 = (nC_st1_b94_c1 == 0) ? nS_st1_b95_c0 : nS_st1_b95_c1;
  assign nS_st2_b96_c1 = nS_st1_b96_c1;
  assign nS_st2_b97_c1 = (nC_st1_b96_c1 == 0) ? nS_st1_b97_c0 : nS_st1_b97_c1;
  assign nS_st2_b98_c1 = nS_st1_b98_c1;
  assign nS_st2_b99_c1 = (nC_st1_b98_c1 == 0) ? nS_st1_b99_c0 : nS_st1_b99_c1;
  assign nS_st2_b100_c1 = nS_st1_b100_c1;
  assign nS_st2_b101_c1 = (nC_st1_b100_c1 == 0) ? nS_st1_b101_c0 : nS_st1_b101_c1;
  assign nS_st2_b102_c1 = nS_st1_b102_c1;
  assign nS_st2_b103_c1 = (nC_st1_b102_c1 == 0) ? nS_st1_b103_c0 : nS_st1_b103_c1;
  assign nS_st2_b104_c1 = nS_st1_b104_c1;
  assign nS_st2_b105_c1 = (nC_st1_b104_c1 == 0) ? nS_st1_b105_c0 : nS_st1_b105_c1;
  assign nS_st2_b106_c1 = nS_st1_b106_c1;
  assign nS_st2_b107_c1 = (nC_st1_b106_c1 == 0) ? nS_st1_b107_c0 : nS_st1_b107_c1;
  assign nS_st2_b108_c1 = nS_st1_b108_c1;
  assign nS_st2_b109_c1 = (nC_st1_b108_c1 == 0) ? nS_st1_b109_c0 : nS_st1_b109_c1;
  assign nS_st2_b110_c1 = nS_st1_b110_c1;
  assign nS_st2_b111_c1 = (nC_st1_b110_c1 == 0) ? nS_st1_b111_c0 : nS_st1_b111_c1;
  assign nS_st2_b112_c1 = nS_st1_b112_c1;
  assign nS_st2_b113_c1 = (nC_st1_b112_c1 == 0) ? nS_st1_b113_c0 : nS_st1_b113_c1;
  assign nS_st2_b114_c1 = nS_st1_b114_c1;
  assign nS_st2_b115_c1 = (nC_st1_b114_c1 == 0) ? nS_st1_b115_c0 : nS_st1_b115_c1;
  assign nS_st2_b116_c1 = nS_st1_b116_c1;
  assign nS_st2_b117_c1 = (nC_st1_b116_c1 == 0) ? nS_st1_b117_c0 : nS_st1_b117_c1;
  assign nS_st2_b118_c1 = nS_st1_b118_c1;
  assign nS_st2_b119_c1 = (nC_st1_b118_c1 == 0) ? nS_st1_b119_c0 : nS_st1_b119_c1;
  assign nS_st2_b120_c1 = nS_st1_b120_c1;
  assign nS_st2_b121_c1 = (nC_st1_b120_c1 == 0) ? nS_st1_b121_c0 : nS_st1_b121_c1;
  assign nS_st2_b122_c1 = nS_st1_b122_c1;
  assign nS_st2_b123_c1 = (nC_st1_b122_c1 == 0) ? nS_st1_b123_c0 : nS_st1_b123_c1;
  assign nS_st2_b124_c1 = nS_st1_b124_c1;
  assign nS_st2_b125_c1 = (nC_st1_b124_c1 == 0) ? nS_st1_b125_c0 : nS_st1_b125_c1;
  assign nS_st2_b126_c1 = nS_st1_b126_c1;
  assign nS_st2_b127_c1 = (nC_st1_b126_c1 == 0) ? nS_st1_b127_c0 : nS_st1_b127_c1;
  assign nC_st2_b1_c0 = (nC_st1_b0_c0 == 0) ? nC_st1_b1_c0 : nC_st1_b1_c1;
  assign nC_st2_b3_c0 = (nC_st1_b2_c0 == 0) ? nC_st1_b3_c0 : nC_st1_b3_c1;
  assign nC_st2_b5_c0 = (nC_st1_b4_c0 == 0) ? nC_st1_b5_c0 : nC_st1_b5_c1;
  assign nC_st2_b7_c0 = (nC_st1_b6_c0 == 0) ? nC_st1_b7_c0 : nC_st1_b7_c1;
  assign nC_st2_b9_c0 = (nC_st1_b8_c0 == 0) ? nC_st1_b9_c0 : nC_st1_b9_c1;
  assign nC_st2_b11_c0 = (nC_st1_b10_c0 == 0) ? nC_st1_b11_c0 : nC_st1_b11_c1;
  assign nC_st2_b13_c0 = (nC_st1_b12_c0 == 0) ? nC_st1_b13_c0 : nC_st1_b13_c1;
  assign nC_st2_b15_c0 = (nC_st1_b14_c0 == 0) ? nC_st1_b15_c0 : nC_st1_b15_c1;
  assign nC_st2_b17_c0 = (nC_st1_b16_c0 == 0) ? nC_st1_b17_c0 : nC_st1_b17_c1;
  assign nC_st2_b19_c0 = (nC_st1_b18_c0 == 0) ? nC_st1_b19_c0 : nC_st1_b19_c1;
  assign nC_st2_b21_c0 = (nC_st1_b20_c0 == 0) ? nC_st1_b21_c0 : nC_st1_b21_c1;
  assign nC_st2_b23_c0 = (nC_st1_b22_c0 == 0) ? nC_st1_b23_c0 : nC_st1_b23_c1;
  assign nC_st2_b25_c0 = (nC_st1_b24_c0 == 0) ? nC_st1_b25_c0 : nC_st1_b25_c1;
  assign nC_st2_b27_c0 = (nC_st1_b26_c0 == 0) ? nC_st1_b27_c0 : nC_st1_b27_c1;
  assign nC_st2_b29_c0 = (nC_st1_b28_c0 == 0) ? nC_st1_b29_c0 : nC_st1_b29_c1;
  assign nC_st2_b31_c0 = (nC_st1_b30_c0 == 0) ? nC_st1_b31_c0 : nC_st1_b31_c1;
  assign nC_st2_b33_c0 = (nC_st1_b32_c0 == 0) ? nC_st1_b33_c0 : nC_st1_b33_c1;
  assign nC_st2_b35_c0 = (nC_st1_b34_c0 == 0) ? nC_st1_b35_c0 : nC_st1_b35_c1;
  assign nC_st2_b37_c0 = (nC_st1_b36_c0 == 0) ? nC_st1_b37_c0 : nC_st1_b37_c1;
  assign nC_st2_b39_c0 = (nC_st1_b38_c0 == 0) ? nC_st1_b39_c0 : nC_st1_b39_c1;
  assign nC_st2_b41_c0 = (nC_st1_b40_c0 == 0) ? nC_st1_b41_c0 : nC_st1_b41_c1;
  assign nC_st2_b43_c0 = (nC_st1_b42_c0 == 0) ? nC_st1_b43_c0 : nC_st1_b43_c1;
  assign nC_st2_b45_c0 = (nC_st1_b44_c0 == 0) ? nC_st1_b45_c0 : nC_st1_b45_c1;
  assign nC_st2_b47_c0 = (nC_st1_b46_c0 == 0) ? nC_st1_b47_c0 : nC_st1_b47_c1;
  assign nC_st2_b49_c0 = (nC_st1_b48_c0 == 0) ? nC_st1_b49_c0 : nC_st1_b49_c1;
  assign nC_st2_b51_c0 = (nC_st1_b50_c0 == 0) ? nC_st1_b51_c0 : nC_st1_b51_c1;
  assign nC_st2_b53_c0 = (nC_st1_b52_c0 == 0) ? nC_st1_b53_c0 : nC_st1_b53_c1;
  assign nC_st2_b55_c0 = (nC_st1_b54_c0 == 0) ? nC_st1_b55_c0 : nC_st1_b55_c1;
  assign nC_st2_b57_c0 = (nC_st1_b56_c0 == 0) ? nC_st1_b57_c0 : nC_st1_b57_c1;
  assign nC_st2_b59_c0 = (nC_st1_b58_c0 == 0) ? nC_st1_b59_c0 : nC_st1_b59_c1;
  assign nC_st2_b61_c0 = (nC_st1_b60_c0 == 0) ? nC_st1_b61_c0 : nC_st1_b61_c1;
  assign nC_st2_b63_c0 = (nC_st1_b62_c0 == 0) ? nC_st1_b63_c0 : nC_st1_b63_c1;
  assign nC_st2_b65_c0 = (nC_st1_b64_c0 == 0) ? nC_st1_b65_c0 : nC_st1_b65_c1;
  assign nC_st2_b67_c0 = (nC_st1_b66_c0 == 0) ? nC_st1_b67_c0 : nC_st1_b67_c1;
  assign nC_st2_b69_c0 = (nC_st1_b68_c0 == 0) ? nC_st1_b69_c0 : nC_st1_b69_c1;
  assign nC_st2_b71_c0 = (nC_st1_b70_c0 == 0) ? nC_st1_b71_c0 : nC_st1_b71_c1;
  assign nC_st2_b73_c0 = (nC_st1_b72_c0 == 0) ? nC_st1_b73_c0 : nC_st1_b73_c1;
  assign nC_st2_b75_c0 = (nC_st1_b74_c0 == 0) ? nC_st1_b75_c0 : nC_st1_b75_c1;
  assign nC_st2_b77_c0 = (nC_st1_b76_c0 == 0) ? nC_st1_b77_c0 : nC_st1_b77_c1;
  assign nC_st2_b79_c0 = (nC_st1_b78_c0 == 0) ? nC_st1_b79_c0 : nC_st1_b79_c1;
  assign nC_st2_b81_c0 = (nC_st1_b80_c0 == 0) ? nC_st1_b81_c0 : nC_st1_b81_c1;
  assign nC_st2_b83_c0 = (nC_st1_b82_c0 == 0) ? nC_st1_b83_c0 : nC_st1_b83_c1;
  assign nC_st2_b85_c0 = (nC_st1_b84_c0 == 0) ? nC_st1_b85_c0 : nC_st1_b85_c1;
  assign nC_st2_b87_c0 = (nC_st1_b86_c0 == 0) ? nC_st1_b87_c0 : nC_st1_b87_c1;
  assign nC_st2_b89_c0 = (nC_st1_b88_c0 == 0) ? nC_st1_b89_c0 : nC_st1_b89_c1;
  assign nC_st2_b91_c0 = (nC_st1_b90_c0 == 0) ? nC_st1_b91_c0 : nC_st1_b91_c1;
  assign nC_st2_b93_c0 = (nC_st1_b92_c0 == 0) ? nC_st1_b93_c0 : nC_st1_b93_c1;
  assign nC_st2_b95_c0 = (nC_st1_b94_c0 == 0) ? nC_st1_b95_c0 : nC_st1_b95_c1;
  assign nC_st2_b97_c0 = (nC_st1_b96_c0 == 0) ? nC_st1_b97_c0 : nC_st1_b97_c1;
  assign nC_st2_b99_c0 = (nC_st1_b98_c0 == 0) ? nC_st1_b99_c0 : nC_st1_b99_c1;
  assign nC_st2_b101_c0 = (nC_st1_b100_c0 == 0) ? nC_st1_b101_c0 : nC_st1_b101_c1;
  assign nC_st2_b103_c0 = (nC_st1_b102_c0 == 0) ? nC_st1_b103_c0 : nC_st1_b103_c1;
  assign nC_st2_b105_c0 = (nC_st1_b104_c0 == 0) ? nC_st1_b105_c0 : nC_st1_b105_c1;
  assign nC_st2_b107_c0 = (nC_st1_b106_c0 == 0) ? nC_st1_b107_c0 : nC_st1_b107_c1;
  assign nC_st2_b109_c0 = (nC_st1_b108_c0 == 0) ? nC_st1_b109_c0 : nC_st1_b109_c1;
  assign nC_st2_b111_c0 = (nC_st1_b110_c0 == 0) ? nC_st1_b111_c0 : nC_st1_b111_c1;
  assign nC_st2_b113_c0 = (nC_st1_b112_c0 == 0) ? nC_st1_b113_c0 : nC_st1_b113_c1;
  assign nC_st2_b115_c0 = (nC_st1_b114_c0 == 0) ? nC_st1_b115_c0 : nC_st1_b115_c1;
  assign nC_st2_b117_c0 = (nC_st1_b116_c0 == 0) ? nC_st1_b117_c0 : nC_st1_b117_c1;
  assign nC_st2_b119_c0 = (nC_st1_b118_c0 == 0) ? nC_st1_b119_c0 : nC_st1_b119_c1;
  assign nC_st2_b121_c0 = (nC_st1_b120_c0 == 0) ? nC_st1_b121_c0 : nC_st1_b121_c1;
  assign nC_st2_b123_c0 = (nC_st1_b122_c0 == 0) ? nC_st1_b123_c0 : nC_st1_b123_c1;
  assign nC_st2_b125_c0 = (nC_st1_b124_c0 == 0) ? nC_st1_b125_c0 : nC_st1_b125_c1;
  assign nC_st2_b127_c0 = (nC_st1_b126_c0 == 0) ? nC_st1_b127_c0 : nC_st1_b127_c1;
  assign nC_st2_b1_c1 = (nC_st1_b0_c1 == 0) ? nC_st1_b1_c0 : nC_st1_b1_c1;
  assign nC_st2_b3_c1 = (nC_st1_b2_c1 == 0) ? nC_st1_b3_c0 : nC_st1_b3_c1;
  assign nC_st2_b5_c1 = (nC_st1_b4_c1 == 0) ? nC_st1_b5_c0 : nC_st1_b5_c1;
  assign nC_st2_b7_c1 = (nC_st1_b6_c1 == 0) ? nC_st1_b7_c0 : nC_st1_b7_c1;
  assign nC_st2_b9_c1 = (nC_st1_b8_c1 == 0) ? nC_st1_b9_c0 : nC_st1_b9_c1;
  assign nC_st2_b11_c1 = (nC_st1_b10_c1 == 0) ? nC_st1_b11_c0 : nC_st1_b11_c1;
  assign nC_st2_b13_c1 = (nC_st1_b12_c1 == 0) ? nC_st1_b13_c0 : nC_st1_b13_c1;
  assign nC_st2_b15_c1 = (nC_st1_b14_c1 == 0) ? nC_st1_b15_c0 : nC_st1_b15_c1;
  assign nC_st2_b17_c1 = (nC_st1_b16_c1 == 0) ? nC_st1_b17_c0 : nC_st1_b17_c1;
  assign nC_st2_b19_c1 = (nC_st1_b18_c1 == 0) ? nC_st1_b19_c0 : nC_st1_b19_c1;
  assign nC_st2_b21_c1 = (nC_st1_b20_c1 == 0) ? nC_st1_b21_c0 : nC_st1_b21_c1;
  assign nC_st2_b23_c1 = (nC_st1_b22_c1 == 0) ? nC_st1_b23_c0 : nC_st1_b23_c1;
  assign nC_st2_b25_c1 = (nC_st1_b24_c1 == 0) ? nC_st1_b25_c0 : nC_st1_b25_c1;
  assign nC_st2_b27_c1 = (nC_st1_b26_c1 == 0) ? nC_st1_b27_c0 : nC_st1_b27_c1;
  assign nC_st2_b29_c1 = (nC_st1_b28_c1 == 0) ? nC_st1_b29_c0 : nC_st1_b29_c1;
  assign nC_st2_b31_c1 = (nC_st1_b30_c1 == 0) ? nC_st1_b31_c0 : nC_st1_b31_c1;
  assign nC_st2_b33_c1 = (nC_st1_b32_c1 == 0) ? nC_st1_b33_c0 : nC_st1_b33_c1;
  assign nC_st2_b35_c1 = (nC_st1_b34_c1 == 0) ? nC_st1_b35_c0 : nC_st1_b35_c1;
  assign nC_st2_b37_c1 = (nC_st1_b36_c1 == 0) ? nC_st1_b37_c0 : nC_st1_b37_c1;
  assign nC_st2_b39_c1 = (nC_st1_b38_c1 == 0) ? nC_st1_b39_c0 : nC_st1_b39_c1;
  assign nC_st2_b41_c1 = (nC_st1_b40_c1 == 0) ? nC_st1_b41_c0 : nC_st1_b41_c1;
  assign nC_st2_b43_c1 = (nC_st1_b42_c1 == 0) ? nC_st1_b43_c0 : nC_st1_b43_c1;
  assign nC_st2_b45_c1 = (nC_st1_b44_c1 == 0) ? nC_st1_b45_c0 : nC_st1_b45_c1;
  assign nC_st2_b47_c1 = (nC_st1_b46_c1 == 0) ? nC_st1_b47_c0 : nC_st1_b47_c1;
  assign nC_st2_b49_c1 = (nC_st1_b48_c1 == 0) ? nC_st1_b49_c0 : nC_st1_b49_c1;
  assign nC_st2_b51_c1 = (nC_st1_b50_c1 == 0) ? nC_st1_b51_c0 : nC_st1_b51_c1;
  assign nC_st2_b53_c1 = (nC_st1_b52_c1 == 0) ? nC_st1_b53_c0 : nC_st1_b53_c1;
  assign nC_st2_b55_c1 = (nC_st1_b54_c1 == 0) ? nC_st1_b55_c0 : nC_st1_b55_c1;
  assign nC_st2_b57_c1 = (nC_st1_b56_c1 == 0) ? nC_st1_b57_c0 : nC_st1_b57_c1;
  assign nC_st2_b59_c1 = (nC_st1_b58_c1 == 0) ? nC_st1_b59_c0 : nC_st1_b59_c1;
  assign nC_st2_b61_c1 = (nC_st1_b60_c1 == 0) ? nC_st1_b61_c0 : nC_st1_b61_c1;
  assign nC_st2_b63_c1 = (nC_st1_b62_c1 == 0) ? nC_st1_b63_c0 : nC_st1_b63_c1;
  assign nC_st2_b65_c1 = (nC_st1_b64_c1 == 0) ? nC_st1_b65_c0 : nC_st1_b65_c1;
  assign nC_st2_b67_c1 = (nC_st1_b66_c1 == 0) ? nC_st1_b67_c0 : nC_st1_b67_c1;
  assign nC_st2_b69_c1 = (nC_st1_b68_c1 == 0) ? nC_st1_b69_c0 : nC_st1_b69_c1;
  assign nC_st2_b71_c1 = (nC_st1_b70_c1 == 0) ? nC_st1_b71_c0 : nC_st1_b71_c1;
  assign nC_st2_b73_c1 = (nC_st1_b72_c1 == 0) ? nC_st1_b73_c0 : nC_st1_b73_c1;
  assign nC_st2_b75_c1 = (nC_st1_b74_c1 == 0) ? nC_st1_b75_c0 : nC_st1_b75_c1;
  assign nC_st2_b77_c1 = (nC_st1_b76_c1 == 0) ? nC_st1_b77_c0 : nC_st1_b77_c1;
  assign nC_st2_b79_c1 = (nC_st1_b78_c1 == 0) ? nC_st1_b79_c0 : nC_st1_b79_c1;
  assign nC_st2_b81_c1 = (nC_st1_b80_c1 == 0) ? nC_st1_b81_c0 : nC_st1_b81_c1;
  assign nC_st2_b83_c1 = (nC_st1_b82_c1 == 0) ? nC_st1_b83_c0 : nC_st1_b83_c1;
  assign nC_st2_b85_c1 = (nC_st1_b84_c1 == 0) ? nC_st1_b85_c0 : nC_st1_b85_c1;
  assign nC_st2_b87_c1 = (nC_st1_b86_c1 == 0) ? nC_st1_b87_c0 : nC_st1_b87_c1;
  assign nC_st2_b89_c1 = (nC_st1_b88_c1 == 0) ? nC_st1_b89_c0 : nC_st1_b89_c1;
  assign nC_st2_b91_c1 = (nC_st1_b90_c1 == 0) ? nC_st1_b91_c0 : nC_st1_b91_c1;
  assign nC_st2_b93_c1 = (nC_st1_b92_c1 == 0) ? nC_st1_b93_c0 : nC_st1_b93_c1;
  assign nC_st2_b95_c1 = (nC_st1_b94_c1 == 0) ? nC_st1_b95_c0 : nC_st1_b95_c1;
  assign nC_st2_b97_c1 = (nC_st1_b96_c1 == 0) ? nC_st1_b97_c0 : nC_st1_b97_c1;
  assign nC_st2_b99_c1 = (nC_st1_b98_c1 == 0) ? nC_st1_b99_c0 : nC_st1_b99_c1;
  assign nC_st2_b101_c1 = (nC_st1_b100_c1 == 0) ? nC_st1_b101_c0 : nC_st1_b101_c1;
  assign nC_st2_b103_c1 = (nC_st1_b102_c1 == 0) ? nC_st1_b103_c0 : nC_st1_b103_c1;
  assign nC_st2_b105_c1 = (nC_st1_b104_c1 == 0) ? nC_st1_b105_c0 : nC_st1_b105_c1;
  assign nC_st2_b107_c1 = (nC_st1_b106_c1 == 0) ? nC_st1_b107_c0 : nC_st1_b107_c1;
  assign nC_st2_b109_c1 = (nC_st1_b108_c1 == 0) ? nC_st1_b109_c0 : nC_st1_b109_c1;
  assign nC_st2_b111_c1 = (nC_st1_b110_c1 == 0) ? nC_st1_b111_c0 : nC_st1_b111_c1;
  assign nC_st2_b113_c1 = (nC_st1_b112_c1 == 0) ? nC_st1_b113_c0 : nC_st1_b113_c1;
  assign nC_st2_b115_c1 = (nC_st1_b114_c1 == 0) ? nC_st1_b115_c0 : nC_st1_b115_c1;
  assign nC_st2_b117_c1 = (nC_st1_b116_c1 == 0) ? nC_st1_b117_c0 : nC_st1_b117_c1;
  assign nC_st2_b119_c1 = (nC_st1_b118_c1 == 0) ? nC_st1_b119_c0 : nC_st1_b119_c1;
  assign nC_st2_b121_c1 = (nC_st1_b120_c1 == 0) ? nC_st1_b121_c0 : nC_st1_b121_c1;
  assign nC_st2_b123_c1 = (nC_st1_b122_c1 == 0) ? nC_st1_b123_c0 : nC_st1_b123_c1;
  assign nC_st2_b125_c1 = (nC_st1_b124_c1 == 0) ? nC_st1_b125_c0 : nC_st1_b125_c1;
  assign nC_st2_b127_c1 = (nC_st1_b126_c1 == 0) ? nC_st1_b127_c0 : nC_st1_b127_c1;

  assign nS_st3_b0_c0 = nS_st2_b0_c0;
  assign nS_st3_b1_c0 = nS_st2_b1_c0;
  assign nS_st3_b2_c0 = (nC_st2_b1_c0 == 0) ? nS_st2_b2_c0 : nS_st2_b2_c1;
  assign nS_st3_b3_c0 = (nC_st2_b1_c0 == 0) ? nS_st2_b3_c0 : nS_st2_b3_c1;
  assign nS_st3_b4_c0 = nS_st2_b4_c0;
  assign nS_st3_b5_c0 = nS_st2_b5_c0;
  assign nS_st3_b6_c0 = (nC_st2_b5_c0 == 0) ? nS_st2_b6_c0 : nS_st2_b6_c1;
  assign nS_st3_b7_c0 = (nC_st2_b5_c0 == 0) ? nS_st2_b7_c0 : nS_st2_b7_c1;
  assign nS_st3_b8_c0 = nS_st2_b8_c0;
  assign nS_st3_b9_c0 = nS_st2_b9_c0;
  assign nS_st3_b10_c0 = (nC_st2_b9_c0 == 0) ? nS_st2_b10_c0 : nS_st2_b10_c1;
  assign nS_st3_b11_c0 = (nC_st2_b9_c0 == 0) ? nS_st2_b11_c0 : nS_st2_b11_c1;
  assign nS_st3_b12_c0 = nS_st2_b12_c0;
  assign nS_st3_b13_c0 = nS_st2_b13_c0;
  assign nS_st3_b14_c0 = (nC_st2_b13_c0 == 0) ? nS_st2_b14_c0 : nS_st2_b14_c1;
  assign nS_st3_b15_c0 = (nC_st2_b13_c0 == 0) ? nS_st2_b15_c0 : nS_st2_b15_c1;
  assign nS_st3_b16_c0 = nS_st2_b16_c0;
  assign nS_st3_b17_c0 = nS_st2_b17_c0;
  assign nS_st3_b18_c0 = (nC_st2_b17_c0 == 0) ? nS_st2_b18_c0 : nS_st2_b18_c1;
  assign nS_st3_b19_c0 = (nC_st2_b17_c0 == 0) ? nS_st2_b19_c0 : nS_st2_b19_c1;
  assign nS_st3_b20_c0 = nS_st2_b20_c0;
  assign nS_st3_b21_c0 = nS_st2_b21_c0;
  assign nS_st3_b22_c0 = (nC_st2_b21_c0 == 0) ? nS_st2_b22_c0 : nS_st2_b22_c1;
  assign nS_st3_b23_c0 = (nC_st2_b21_c0 == 0) ? nS_st2_b23_c0 : nS_st2_b23_c1;
  assign nS_st3_b24_c0 = nS_st2_b24_c0;
  assign nS_st3_b25_c0 = nS_st2_b25_c0;
  assign nS_st3_b26_c0 = (nC_st2_b25_c0 == 0) ? nS_st2_b26_c0 : nS_st2_b26_c1;
  assign nS_st3_b27_c0 = (nC_st2_b25_c0 == 0) ? nS_st2_b27_c0 : nS_st2_b27_c1;
  assign nS_st3_b28_c0 = nS_st2_b28_c0;
  assign nS_st3_b29_c0 = nS_st2_b29_c0;
  assign nS_st3_b30_c0 = (nC_st2_b29_c0 == 0) ? nS_st2_b30_c0 : nS_st2_b30_c1;
  assign nS_st3_b31_c0 = (nC_st2_b29_c0 == 0) ? nS_st2_b31_c0 : nS_st2_b31_c1;
  assign nS_st3_b32_c0 = nS_st2_b32_c0;
  assign nS_st3_b33_c0 = nS_st2_b33_c0;
  assign nS_st3_b34_c0 = (nC_st2_b33_c0 == 0) ? nS_st2_b34_c0 : nS_st2_b34_c1;
  assign nS_st3_b35_c0 = (nC_st2_b33_c0 == 0) ? nS_st2_b35_c0 : nS_st2_b35_c1;
  assign nS_st3_b36_c0 = nS_st2_b36_c0;
  assign nS_st3_b37_c0 = nS_st2_b37_c0;
  assign nS_st3_b38_c0 = (nC_st2_b37_c0 == 0) ? nS_st2_b38_c0 : nS_st2_b38_c1;
  assign nS_st3_b39_c0 = (nC_st2_b37_c0 == 0) ? nS_st2_b39_c0 : nS_st2_b39_c1;
  assign nS_st3_b40_c0 = nS_st2_b40_c0;
  assign nS_st3_b41_c0 = nS_st2_b41_c0;
  assign nS_st3_b42_c0 = (nC_st2_b41_c0 == 0) ? nS_st2_b42_c0 : nS_st2_b42_c1;
  assign nS_st3_b43_c0 = (nC_st2_b41_c0 == 0) ? nS_st2_b43_c0 : nS_st2_b43_c1;
  assign nS_st3_b44_c0 = nS_st2_b44_c0;
  assign nS_st3_b45_c0 = nS_st2_b45_c0;
  assign nS_st3_b46_c0 = (nC_st2_b45_c0 == 0) ? nS_st2_b46_c0 : nS_st2_b46_c1;
  assign nS_st3_b47_c0 = (nC_st2_b45_c0 == 0) ? nS_st2_b47_c0 : nS_st2_b47_c1;
  assign nS_st3_b48_c0 = nS_st2_b48_c0;
  assign nS_st3_b49_c0 = nS_st2_b49_c0;
  assign nS_st3_b50_c0 = (nC_st2_b49_c0 == 0) ? nS_st2_b50_c0 : nS_st2_b50_c1;
  assign nS_st3_b51_c0 = (nC_st2_b49_c0 == 0) ? nS_st2_b51_c0 : nS_st2_b51_c1;
  assign nS_st3_b52_c0 = nS_st2_b52_c0;
  assign nS_st3_b53_c0 = nS_st2_b53_c0;
  assign nS_st3_b54_c0 = (nC_st2_b53_c0 == 0) ? nS_st2_b54_c0 : nS_st2_b54_c1;
  assign nS_st3_b55_c0 = (nC_st2_b53_c0 == 0) ? nS_st2_b55_c0 : nS_st2_b55_c1;
  assign nS_st3_b56_c0 = nS_st2_b56_c0;
  assign nS_st3_b57_c0 = nS_st2_b57_c0;
  assign nS_st3_b58_c0 = (nC_st2_b57_c0 == 0) ? nS_st2_b58_c0 : nS_st2_b58_c1;
  assign nS_st3_b59_c0 = (nC_st2_b57_c0 == 0) ? nS_st2_b59_c0 : nS_st2_b59_c1;
  assign nS_st3_b60_c0 = nS_st2_b60_c0;
  assign nS_st3_b61_c0 = nS_st2_b61_c0;
  assign nS_st3_b62_c0 = (nC_st2_b61_c0 == 0) ? nS_st2_b62_c0 : nS_st2_b62_c1;
  assign nS_st3_b63_c0 = (nC_st2_b61_c0 == 0) ? nS_st2_b63_c0 : nS_st2_b63_c1;
  assign nS_st3_b64_c0 = nS_st2_b64_c0;
  assign nS_st3_b65_c0 = nS_st2_b65_c0;
  assign nS_st3_b66_c0 = (nC_st2_b65_c0 == 0) ? nS_st2_b66_c0 : nS_st2_b66_c1;
  assign nS_st3_b67_c0 = (nC_st2_b65_c0 == 0) ? nS_st2_b67_c0 : nS_st2_b67_c1;
  assign nS_st3_b68_c0 = nS_st2_b68_c0;
  assign nS_st3_b69_c0 = nS_st2_b69_c0;
  assign nS_st3_b70_c0 = (nC_st2_b69_c0 == 0) ? nS_st2_b70_c0 : nS_st2_b70_c1;
  assign nS_st3_b71_c0 = (nC_st2_b69_c0 == 0) ? nS_st2_b71_c0 : nS_st2_b71_c1;
  assign nS_st3_b72_c0 = nS_st2_b72_c0;
  assign nS_st3_b73_c0 = nS_st2_b73_c0;
  assign nS_st3_b74_c0 = (nC_st2_b73_c0 == 0) ? nS_st2_b74_c0 : nS_st2_b74_c1;
  assign nS_st3_b75_c0 = (nC_st2_b73_c0 == 0) ? nS_st2_b75_c0 : nS_st2_b75_c1;
  assign nS_st3_b76_c0 = nS_st2_b76_c0;
  assign nS_st3_b77_c0 = nS_st2_b77_c0;
  assign nS_st3_b78_c0 = (nC_st2_b77_c0 == 0) ? nS_st2_b78_c0 : nS_st2_b78_c1;
  assign nS_st3_b79_c0 = (nC_st2_b77_c0 == 0) ? nS_st2_b79_c0 : nS_st2_b79_c1;
  assign nS_st3_b80_c0 = nS_st2_b80_c0;
  assign nS_st3_b81_c0 = nS_st2_b81_c0;
  assign nS_st3_b82_c0 = (nC_st2_b81_c0 == 0) ? nS_st2_b82_c0 : nS_st2_b82_c1;
  assign nS_st3_b83_c0 = (nC_st2_b81_c0 == 0) ? nS_st2_b83_c0 : nS_st2_b83_c1;
  assign nS_st3_b84_c0 = nS_st2_b84_c0;
  assign nS_st3_b85_c0 = nS_st2_b85_c0;
  assign nS_st3_b86_c0 = (nC_st2_b85_c0 == 0) ? nS_st2_b86_c0 : nS_st2_b86_c1;
  assign nS_st3_b87_c0 = (nC_st2_b85_c0 == 0) ? nS_st2_b87_c0 : nS_st2_b87_c1;
  assign nS_st3_b88_c0 = nS_st2_b88_c0;
  assign nS_st3_b89_c0 = nS_st2_b89_c0;
  assign nS_st3_b90_c0 = (nC_st2_b89_c0 == 0) ? nS_st2_b90_c0 : nS_st2_b90_c1;
  assign nS_st3_b91_c0 = (nC_st2_b89_c0 == 0) ? nS_st2_b91_c0 : nS_st2_b91_c1;
  assign nS_st3_b92_c0 = nS_st2_b92_c0;
  assign nS_st3_b93_c0 = nS_st2_b93_c0;
  assign nS_st3_b94_c0 = (nC_st2_b93_c0 == 0) ? nS_st2_b94_c0 : nS_st2_b94_c1;
  assign nS_st3_b95_c0 = (nC_st2_b93_c0 == 0) ? nS_st2_b95_c0 : nS_st2_b95_c1;
  assign nS_st3_b96_c0 = nS_st2_b96_c0;
  assign nS_st3_b97_c0 = nS_st2_b97_c0;
  assign nS_st3_b98_c0 = (nC_st2_b97_c0 == 0) ? nS_st2_b98_c0 : nS_st2_b98_c1;
  assign nS_st3_b99_c0 = (nC_st2_b97_c0 == 0) ? nS_st2_b99_c0 : nS_st2_b99_c1;
  assign nS_st3_b100_c0 = nS_st2_b100_c0;
  assign nS_st3_b101_c0 = nS_st2_b101_c0;
  assign nS_st3_b102_c0 = (nC_st2_b101_c0 == 0) ? nS_st2_b102_c0 : nS_st2_b102_c1;
  assign nS_st3_b103_c0 = (nC_st2_b101_c0 == 0) ? nS_st2_b103_c0 : nS_st2_b103_c1;
  assign nS_st3_b104_c0 = nS_st2_b104_c0;
  assign nS_st3_b105_c0 = nS_st2_b105_c0;
  assign nS_st3_b106_c0 = (nC_st2_b105_c0 == 0) ? nS_st2_b106_c0 : nS_st2_b106_c1;
  assign nS_st3_b107_c0 = (nC_st2_b105_c0 == 0) ? nS_st2_b107_c0 : nS_st2_b107_c1;
  assign nS_st3_b108_c0 = nS_st2_b108_c0;
  assign nS_st3_b109_c0 = nS_st2_b109_c0;
  assign nS_st3_b110_c0 = (nC_st2_b109_c0 == 0) ? nS_st2_b110_c0 : nS_st2_b110_c1;
  assign nS_st3_b111_c0 = (nC_st2_b109_c0 == 0) ? nS_st2_b111_c0 : nS_st2_b111_c1;
  assign nS_st3_b112_c0 = nS_st2_b112_c0;
  assign nS_st3_b113_c0 = nS_st2_b113_c0;
  assign nS_st3_b114_c0 = (nC_st2_b113_c0 == 0) ? nS_st2_b114_c0 : nS_st2_b114_c1;
  assign nS_st3_b115_c0 = (nC_st2_b113_c0 == 0) ? nS_st2_b115_c0 : nS_st2_b115_c1;
  assign nS_st3_b116_c0 = nS_st2_b116_c0;
  assign nS_st3_b117_c0 = nS_st2_b117_c0;
  assign nS_st3_b118_c0 = (nC_st2_b117_c0 == 0) ? nS_st2_b118_c0 : nS_st2_b118_c1;
  assign nS_st3_b119_c0 = (nC_st2_b117_c0 == 0) ? nS_st2_b119_c0 : nS_st2_b119_c1;
  assign nS_st3_b120_c0 = nS_st2_b120_c0;
  assign nS_st3_b121_c0 = nS_st2_b121_c0;
  assign nS_st3_b122_c0 = (nC_st2_b121_c0 == 0) ? nS_st2_b122_c0 : nS_st2_b122_c1;
  assign nS_st3_b123_c0 = (nC_st2_b121_c0 == 0) ? nS_st2_b123_c0 : nS_st2_b123_c1;
  assign nS_st3_b124_c0 = nS_st2_b124_c0;
  assign nS_st3_b125_c0 = nS_st2_b125_c0;
  assign nS_st3_b126_c0 = (nC_st2_b125_c0 == 0) ? nS_st2_b126_c0 : nS_st2_b126_c1;
  assign nS_st3_b127_c0 = (nC_st2_b125_c0 == 0) ? nS_st2_b127_c0 : nS_st2_b127_c1;
  assign nS_st3_b0_c1 = nS_st2_b0_c1;
  assign nS_st3_b1_c1 = nS_st2_b1_c1;
  assign nS_st3_b2_c1 = (nC_st2_b1_c1 == 0) ? nS_st2_b2_c0 : nS_st2_b2_c1;
  assign nS_st3_b3_c1 = (nC_st2_b1_c1 == 0) ? nS_st2_b3_c0 : nS_st2_b3_c1;
  assign nS_st3_b4_c1 = nS_st2_b4_c1;
  assign nS_st3_b5_c1 = nS_st2_b5_c1;
  assign nS_st3_b6_c1 = (nC_st2_b5_c1 == 0) ? nS_st2_b6_c0 : nS_st2_b6_c1;
  assign nS_st3_b7_c1 = (nC_st2_b5_c1 == 0) ? nS_st2_b7_c0 : nS_st2_b7_c1;
  assign nS_st3_b8_c1 = nS_st2_b8_c1;
  assign nS_st3_b9_c1 = nS_st2_b9_c1;
  assign nS_st3_b10_c1 = (nC_st2_b9_c1 == 0) ? nS_st2_b10_c0 : nS_st2_b10_c1;
  assign nS_st3_b11_c1 = (nC_st2_b9_c1 == 0) ? nS_st2_b11_c0 : nS_st2_b11_c1;
  assign nS_st3_b12_c1 = nS_st2_b12_c1;
  assign nS_st3_b13_c1 = nS_st2_b13_c1;
  assign nS_st3_b14_c1 = (nC_st2_b13_c1 == 0) ? nS_st2_b14_c0 : nS_st2_b14_c1;
  assign nS_st3_b15_c1 = (nC_st2_b13_c1 == 0) ? nS_st2_b15_c0 : nS_st2_b15_c1;
  assign nS_st3_b16_c1 = nS_st2_b16_c1;
  assign nS_st3_b17_c1 = nS_st2_b17_c1;
  assign nS_st3_b18_c1 = (nC_st2_b17_c1 == 0) ? nS_st2_b18_c0 : nS_st2_b18_c1;
  assign nS_st3_b19_c1 = (nC_st2_b17_c1 == 0) ? nS_st2_b19_c0 : nS_st2_b19_c1;
  assign nS_st3_b20_c1 = nS_st2_b20_c1;
  assign nS_st3_b21_c1 = nS_st2_b21_c1;
  assign nS_st3_b22_c1 = (nC_st2_b21_c1 == 0) ? nS_st2_b22_c0 : nS_st2_b22_c1;
  assign nS_st3_b23_c1 = (nC_st2_b21_c1 == 0) ? nS_st2_b23_c0 : nS_st2_b23_c1;
  assign nS_st3_b24_c1 = nS_st2_b24_c1;
  assign nS_st3_b25_c1 = nS_st2_b25_c1;
  assign nS_st3_b26_c1 = (nC_st2_b25_c1 == 0) ? nS_st2_b26_c0 : nS_st2_b26_c1;
  assign nS_st3_b27_c1 = (nC_st2_b25_c1 == 0) ? nS_st2_b27_c0 : nS_st2_b27_c1;
  assign nS_st3_b28_c1 = nS_st2_b28_c1;
  assign nS_st3_b29_c1 = nS_st2_b29_c1;
  assign nS_st3_b30_c1 = (nC_st2_b29_c1 == 0) ? nS_st2_b30_c0 : nS_st2_b30_c1;
  assign nS_st3_b31_c1 = (nC_st2_b29_c1 == 0) ? nS_st2_b31_c0 : nS_st2_b31_c1;
  assign nS_st3_b32_c1 = nS_st2_b32_c1;
  assign nS_st3_b33_c1 = nS_st2_b33_c1;
  assign nS_st3_b34_c1 = (nC_st2_b33_c1 == 0) ? nS_st2_b34_c0 : nS_st2_b34_c1;
  assign nS_st3_b35_c1 = (nC_st2_b33_c1 == 0) ? nS_st2_b35_c0 : nS_st2_b35_c1;
  assign nS_st3_b36_c1 = nS_st2_b36_c1;
  assign nS_st3_b37_c1 = nS_st2_b37_c1;
  assign nS_st3_b38_c1 = (nC_st2_b37_c1 == 0) ? nS_st2_b38_c0 : nS_st2_b38_c1;
  assign nS_st3_b39_c1 = (nC_st2_b37_c1 == 0) ? nS_st2_b39_c0 : nS_st2_b39_c1;
  assign nS_st3_b40_c1 = nS_st2_b40_c1;
  assign nS_st3_b41_c1 = nS_st2_b41_c1;
  assign nS_st3_b42_c1 = (nC_st2_b41_c1 == 0) ? nS_st2_b42_c0 : nS_st2_b42_c1;
  assign nS_st3_b43_c1 = (nC_st2_b41_c1 == 0) ? nS_st2_b43_c0 : nS_st2_b43_c1;
  assign nS_st3_b44_c1 = nS_st2_b44_c1;
  assign nS_st3_b45_c1 = nS_st2_b45_c1;
  assign nS_st3_b46_c1 = (nC_st2_b45_c1 == 0) ? nS_st2_b46_c0 : nS_st2_b46_c1;
  assign nS_st3_b47_c1 = (nC_st2_b45_c1 == 0) ? nS_st2_b47_c0 : nS_st2_b47_c1;
  assign nS_st3_b48_c1 = nS_st2_b48_c1;
  assign nS_st3_b49_c1 = nS_st2_b49_c1;
  assign nS_st3_b50_c1 = (nC_st2_b49_c1 == 0) ? nS_st2_b50_c0 : nS_st2_b50_c1;
  assign nS_st3_b51_c1 = (nC_st2_b49_c1 == 0) ? nS_st2_b51_c0 : nS_st2_b51_c1;
  assign nS_st3_b52_c1 = nS_st2_b52_c1;
  assign nS_st3_b53_c1 = nS_st2_b53_c1;
  assign nS_st3_b54_c1 = (nC_st2_b53_c1 == 0) ? nS_st2_b54_c0 : nS_st2_b54_c1;
  assign nS_st3_b55_c1 = (nC_st2_b53_c1 == 0) ? nS_st2_b55_c0 : nS_st2_b55_c1;
  assign nS_st3_b56_c1 = nS_st2_b56_c1;
  assign nS_st3_b57_c1 = nS_st2_b57_c1;
  assign nS_st3_b58_c1 = (nC_st2_b57_c1 == 0) ? nS_st2_b58_c0 : nS_st2_b58_c1;
  assign nS_st3_b59_c1 = (nC_st2_b57_c1 == 0) ? nS_st2_b59_c0 : nS_st2_b59_c1;
  assign nS_st3_b60_c1 = nS_st2_b60_c1;
  assign nS_st3_b61_c1 = nS_st2_b61_c1;
  assign nS_st3_b62_c1 = (nC_st2_b61_c1 == 0) ? nS_st2_b62_c0 : nS_st2_b62_c1;
  assign nS_st3_b63_c1 = (nC_st2_b61_c1 == 0) ? nS_st2_b63_c0 : nS_st2_b63_c1;
  assign nS_st3_b64_c1 = nS_st2_b64_c1;
  assign nS_st3_b65_c1 = nS_st2_b65_c1;
  assign nS_st3_b66_c1 = (nC_st2_b65_c1 == 0) ? nS_st2_b66_c0 : nS_st2_b66_c1;
  assign nS_st3_b67_c1 = (nC_st2_b65_c1 == 0) ? nS_st2_b67_c0 : nS_st2_b67_c1;
  assign nS_st3_b68_c1 = nS_st2_b68_c1;
  assign nS_st3_b69_c1 = nS_st2_b69_c1;
  assign nS_st3_b70_c1 = (nC_st2_b69_c1 == 0) ? nS_st2_b70_c0 : nS_st2_b70_c1;
  assign nS_st3_b71_c1 = (nC_st2_b69_c1 == 0) ? nS_st2_b71_c0 : nS_st2_b71_c1;
  assign nS_st3_b72_c1 = nS_st2_b72_c1;
  assign nS_st3_b73_c1 = nS_st2_b73_c1;
  assign nS_st3_b74_c1 = (nC_st2_b73_c1 == 0) ? nS_st2_b74_c0 : nS_st2_b74_c1;
  assign nS_st3_b75_c1 = (nC_st2_b73_c1 == 0) ? nS_st2_b75_c0 : nS_st2_b75_c1;
  assign nS_st3_b76_c1 = nS_st2_b76_c1;
  assign nS_st3_b77_c1 = nS_st2_b77_c1;
  assign nS_st3_b78_c1 = (nC_st2_b77_c1 == 0) ? nS_st2_b78_c0 : nS_st2_b78_c1;
  assign nS_st3_b79_c1 = (nC_st2_b77_c1 == 0) ? nS_st2_b79_c0 : nS_st2_b79_c1;
  assign nS_st3_b80_c1 = nS_st2_b80_c1;
  assign nS_st3_b81_c1 = nS_st2_b81_c1;
  assign nS_st3_b82_c1 = (nC_st2_b81_c1 == 0) ? nS_st2_b82_c0 : nS_st2_b82_c1;
  assign nS_st3_b83_c1 = (nC_st2_b81_c1 == 0) ? nS_st2_b83_c0 : nS_st2_b83_c1;
  assign nS_st3_b84_c1 = nS_st2_b84_c1;
  assign nS_st3_b85_c1 = nS_st2_b85_c1;
  assign nS_st3_b86_c1 = (nC_st2_b85_c1 == 0) ? nS_st2_b86_c0 : nS_st2_b86_c1;
  assign nS_st3_b87_c1 = (nC_st2_b85_c1 == 0) ? nS_st2_b87_c0 : nS_st2_b87_c1;
  assign nS_st3_b88_c1 = nS_st2_b88_c1;
  assign nS_st3_b89_c1 = nS_st2_b89_c1;
  assign nS_st3_b90_c1 = (nC_st2_b89_c1 == 0) ? nS_st2_b90_c0 : nS_st2_b90_c1;
  assign nS_st3_b91_c1 = (nC_st2_b89_c1 == 0) ? nS_st2_b91_c0 : nS_st2_b91_c1;
  assign nS_st3_b92_c1 = nS_st2_b92_c1;
  assign nS_st3_b93_c1 = nS_st2_b93_c1;
  assign nS_st3_b94_c1 = (nC_st2_b93_c1 == 0) ? nS_st2_b94_c0 : nS_st2_b94_c1;
  assign nS_st3_b95_c1 = (nC_st2_b93_c1 == 0) ? nS_st2_b95_c0 : nS_st2_b95_c1;
  assign nS_st3_b96_c1 = nS_st2_b96_c1;
  assign nS_st3_b97_c1 = nS_st2_b97_c1;
  assign nS_st3_b98_c1 = (nC_st2_b97_c1 == 0) ? nS_st2_b98_c0 : nS_st2_b98_c1;
  assign nS_st3_b99_c1 = (nC_st2_b97_c1 == 0) ? nS_st2_b99_c0 : nS_st2_b99_c1;
  assign nS_st3_b100_c1 = nS_st2_b100_c1;
  assign nS_st3_b101_c1 = nS_st2_b101_c1;
  assign nS_st3_b102_c1 = (nC_st2_b101_c1 == 0) ? nS_st2_b102_c0 : nS_st2_b102_c1;
  assign nS_st3_b103_c1 = (nC_st2_b101_c1 == 0) ? nS_st2_b103_c0 : nS_st2_b103_c1;
  assign nS_st3_b104_c1 = nS_st2_b104_c1;
  assign nS_st3_b105_c1 = nS_st2_b105_c1;
  assign nS_st3_b106_c1 = (nC_st2_b105_c1 == 0) ? nS_st2_b106_c0 : nS_st2_b106_c1;
  assign nS_st3_b107_c1 = (nC_st2_b105_c1 == 0) ? nS_st2_b107_c0 : nS_st2_b107_c1;
  assign nS_st3_b108_c1 = nS_st2_b108_c1;
  assign nS_st3_b109_c1 = nS_st2_b109_c1;
  assign nS_st3_b110_c1 = (nC_st2_b109_c1 == 0) ? nS_st2_b110_c0 : nS_st2_b110_c1;
  assign nS_st3_b111_c1 = (nC_st2_b109_c1 == 0) ? nS_st2_b111_c0 : nS_st2_b111_c1;
  assign nS_st3_b112_c1 = nS_st2_b112_c1;
  assign nS_st3_b113_c1 = nS_st2_b113_c1;
  assign nS_st3_b114_c1 = (nC_st2_b113_c1 == 0) ? nS_st2_b114_c0 : nS_st2_b114_c1;
  assign nS_st3_b115_c1 = (nC_st2_b113_c1 == 0) ? nS_st2_b115_c0 : nS_st2_b115_c1;
  assign nS_st3_b116_c1 = nS_st2_b116_c1;
  assign nS_st3_b117_c1 = nS_st2_b117_c1;
  assign nS_st3_b118_c1 = (nC_st2_b117_c1 == 0) ? nS_st2_b118_c0 : nS_st2_b118_c1;
  assign nS_st3_b119_c1 = (nC_st2_b117_c1 == 0) ? nS_st2_b119_c0 : nS_st2_b119_c1;
  assign nS_st3_b120_c1 = nS_st2_b120_c1;
  assign nS_st3_b121_c1 = nS_st2_b121_c1;
  assign nS_st3_b122_c1 = (nC_st2_b121_c1 == 0) ? nS_st2_b122_c0 : nS_st2_b122_c1;
  assign nS_st3_b123_c1 = (nC_st2_b121_c1 == 0) ? nS_st2_b123_c0 : nS_st2_b123_c1;
  assign nS_st3_b124_c1 = nS_st2_b124_c1;
  assign nS_st3_b125_c1 = nS_st2_b125_c1;
  assign nS_st3_b126_c1 = (nC_st2_b125_c1 == 0) ? nS_st2_b126_c0 : nS_st2_b126_c1;
  assign nS_st3_b127_c1 = (nC_st2_b125_c1 == 0) ? nS_st2_b127_c0 : nS_st2_b127_c1;
  assign nC_st3_b3_c0 = (nC_st2_b1_c0 == 0) ? nC_st2_b3_c0 : nC_st2_b3_c1;
  assign nC_st3_b7_c0 = (nC_st2_b5_c0 == 0) ? nC_st2_b7_c0 : nC_st2_b7_c1;
  assign nC_st3_b11_c0 = (nC_st2_b9_c0 == 0) ? nC_st2_b11_c0 : nC_st2_b11_c1;
  assign nC_st3_b15_c0 = (nC_st2_b13_c0 == 0) ? nC_st2_b15_c0 : nC_st2_b15_c1;
  assign nC_st3_b19_c0 = (nC_st2_b17_c0 == 0) ? nC_st2_b19_c0 : nC_st2_b19_c1;
  assign nC_st3_b23_c0 = (nC_st2_b21_c0 == 0) ? nC_st2_b23_c0 : nC_st2_b23_c1;
  assign nC_st3_b27_c0 = (nC_st2_b25_c0 == 0) ? nC_st2_b27_c0 : nC_st2_b27_c1;
  assign nC_st3_b31_c0 = (nC_st2_b29_c0 == 0) ? nC_st2_b31_c0 : nC_st2_b31_c1;
  assign nC_st3_b35_c0 = (nC_st2_b33_c0 == 0) ? nC_st2_b35_c0 : nC_st2_b35_c1;
  assign nC_st3_b39_c0 = (nC_st2_b37_c0 == 0) ? nC_st2_b39_c0 : nC_st2_b39_c1;
  assign nC_st3_b43_c0 = (nC_st2_b41_c0 == 0) ? nC_st2_b43_c0 : nC_st2_b43_c1;
  assign nC_st3_b47_c0 = (nC_st2_b45_c0 == 0) ? nC_st2_b47_c0 : nC_st2_b47_c1;
  assign nC_st3_b51_c0 = (nC_st2_b49_c0 == 0) ? nC_st2_b51_c0 : nC_st2_b51_c1;
  assign nC_st3_b55_c0 = (nC_st2_b53_c0 == 0) ? nC_st2_b55_c0 : nC_st2_b55_c1;
  assign nC_st3_b59_c0 = (nC_st2_b57_c0 == 0) ? nC_st2_b59_c0 : nC_st2_b59_c1;
  assign nC_st3_b63_c0 = (nC_st2_b61_c0 == 0) ? nC_st2_b63_c0 : nC_st2_b63_c1;
  assign nC_st3_b67_c0 = (nC_st2_b65_c0 == 0) ? nC_st2_b67_c0 : nC_st2_b67_c1;
  assign nC_st3_b71_c0 = (nC_st2_b69_c0 == 0) ? nC_st2_b71_c0 : nC_st2_b71_c1;
  assign nC_st3_b75_c0 = (nC_st2_b73_c0 == 0) ? nC_st2_b75_c0 : nC_st2_b75_c1;
  assign nC_st3_b79_c0 = (nC_st2_b77_c0 == 0) ? nC_st2_b79_c0 : nC_st2_b79_c1;
  assign nC_st3_b83_c0 = (nC_st2_b81_c0 == 0) ? nC_st2_b83_c0 : nC_st2_b83_c1;
  assign nC_st3_b87_c0 = (nC_st2_b85_c0 == 0) ? nC_st2_b87_c0 : nC_st2_b87_c1;
  assign nC_st3_b91_c0 = (nC_st2_b89_c0 == 0) ? nC_st2_b91_c0 : nC_st2_b91_c1;
  assign nC_st3_b95_c0 = (nC_st2_b93_c0 == 0) ? nC_st2_b95_c0 : nC_st2_b95_c1;
  assign nC_st3_b99_c0 = (nC_st2_b97_c0 == 0) ? nC_st2_b99_c0 : nC_st2_b99_c1;
  assign nC_st3_b103_c0 = (nC_st2_b101_c0 == 0) ? nC_st2_b103_c0 : nC_st2_b103_c1;
  assign nC_st3_b107_c0 = (nC_st2_b105_c0 == 0) ? nC_st2_b107_c0 : nC_st2_b107_c1;
  assign nC_st3_b111_c0 = (nC_st2_b109_c0 == 0) ? nC_st2_b111_c0 : nC_st2_b111_c1;
  assign nC_st3_b115_c0 = (nC_st2_b113_c0 == 0) ? nC_st2_b115_c0 : nC_st2_b115_c1;
  assign nC_st3_b119_c0 = (nC_st2_b117_c0 == 0) ? nC_st2_b119_c0 : nC_st2_b119_c1;
  assign nC_st3_b123_c0 = (nC_st2_b121_c0 == 0) ? nC_st2_b123_c0 : nC_st2_b123_c1;
  assign nC_st3_b127_c0 = (nC_st2_b125_c0 == 0) ? nC_st2_b127_c0 : nC_st2_b127_c1;
  assign nC_st3_b3_c1 = (nC_st2_b1_c1 == 0) ? nC_st2_b3_c0 : nC_st2_b3_c1;
  assign nC_st3_b7_c1 = (nC_st2_b5_c1 == 0) ? nC_st2_b7_c0 : nC_st2_b7_c1;
  assign nC_st3_b11_c1 = (nC_st2_b9_c1 == 0) ? nC_st2_b11_c0 : nC_st2_b11_c1;
  assign nC_st3_b15_c1 = (nC_st2_b13_c1 == 0) ? nC_st2_b15_c0 : nC_st2_b15_c1;
  assign nC_st3_b19_c1 = (nC_st2_b17_c1 == 0) ? nC_st2_b19_c0 : nC_st2_b19_c1;
  assign nC_st3_b23_c1 = (nC_st2_b21_c1 == 0) ? nC_st2_b23_c0 : nC_st2_b23_c1;
  assign nC_st3_b27_c1 = (nC_st2_b25_c1 == 0) ? nC_st2_b27_c0 : nC_st2_b27_c1;
  assign nC_st3_b31_c1 = (nC_st2_b29_c1 == 0) ? nC_st2_b31_c0 : nC_st2_b31_c1;
  assign nC_st3_b35_c1 = (nC_st2_b33_c1 == 0) ? nC_st2_b35_c0 : nC_st2_b35_c1;
  assign nC_st3_b39_c1 = (nC_st2_b37_c1 == 0) ? nC_st2_b39_c0 : nC_st2_b39_c1;
  assign nC_st3_b43_c1 = (nC_st2_b41_c1 == 0) ? nC_st2_b43_c0 : nC_st2_b43_c1;
  assign nC_st3_b47_c1 = (nC_st2_b45_c1 == 0) ? nC_st2_b47_c0 : nC_st2_b47_c1;
  assign nC_st3_b51_c1 = (nC_st2_b49_c1 == 0) ? nC_st2_b51_c0 : nC_st2_b51_c1;
  assign nC_st3_b55_c1 = (nC_st2_b53_c1 == 0) ? nC_st2_b55_c0 : nC_st2_b55_c1;
  assign nC_st3_b59_c1 = (nC_st2_b57_c1 == 0) ? nC_st2_b59_c0 : nC_st2_b59_c1;
  assign nC_st3_b63_c1 = (nC_st2_b61_c1 == 0) ? nC_st2_b63_c0 : nC_st2_b63_c1;
  assign nC_st3_b67_c1 = (nC_st2_b65_c1 == 0) ? nC_st2_b67_c0 : nC_st2_b67_c1;
  assign nC_st3_b71_c1 = (nC_st2_b69_c1 == 0) ? nC_st2_b71_c0 : nC_st2_b71_c1;
  assign nC_st3_b75_c1 = (nC_st2_b73_c1 == 0) ? nC_st2_b75_c0 : nC_st2_b75_c1;
  assign nC_st3_b79_c1 = (nC_st2_b77_c1 == 0) ? nC_st2_b79_c0 : nC_st2_b79_c1;
  assign nC_st3_b83_c1 = (nC_st2_b81_c1 == 0) ? nC_st2_b83_c0 : nC_st2_b83_c1;
  assign nC_st3_b87_c1 = (nC_st2_b85_c1 == 0) ? nC_st2_b87_c0 : nC_st2_b87_c1;
  assign nC_st3_b91_c1 = (nC_st2_b89_c1 == 0) ? nC_st2_b91_c0 : nC_st2_b91_c1;
  assign nC_st3_b95_c1 = (nC_st2_b93_c1 == 0) ? nC_st2_b95_c0 : nC_st2_b95_c1;
  assign nC_st3_b99_c1 = (nC_st2_b97_c1 == 0) ? nC_st2_b99_c0 : nC_st2_b99_c1;
  assign nC_st3_b103_c1 = (nC_st2_b101_c1 == 0) ? nC_st2_b103_c0 : nC_st2_b103_c1;
  assign nC_st3_b107_c1 = (nC_st2_b105_c1 == 0) ? nC_st2_b107_c0 : nC_st2_b107_c1;
  assign nC_st3_b111_c1 = (nC_st2_b109_c1 == 0) ? nC_st2_b111_c0 : nC_st2_b111_c1;
  assign nC_st3_b115_c1 = (nC_st2_b113_c1 == 0) ? nC_st2_b115_c0 : nC_st2_b115_c1;
  assign nC_st3_b119_c1 = (nC_st2_b117_c1 == 0) ? nC_st2_b119_c0 : nC_st2_b119_c1;
  assign nC_st3_b123_c1 = (nC_st2_b121_c1 == 0) ? nC_st2_b123_c0 : nC_st2_b123_c1;
  assign nC_st3_b127_c1 = (nC_st2_b125_c1 == 0) ? nC_st2_b127_c0 : nC_st2_b127_c1;

  assign nS_st4_b0_c0 = nS_st3_b0_c0;
  assign nS_st4_b1_c0 = nS_st3_b1_c0;
  assign nS_st4_b2_c0 = nS_st3_b2_c0;
  assign nS_st4_b3_c0 = nS_st3_b3_c0;
  assign nS_st4_b4_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b4_c0 : nS_st3_b4_c1;
  assign nS_st4_b5_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b5_c0 : nS_st3_b5_c1;
  assign nS_st4_b6_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b6_c0 : nS_st3_b6_c1;
  assign nS_st4_b7_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b7_c0 : nS_st3_b7_c1;
  assign nS_st4_b8_c0 = nS_st3_b8_c0;
  assign nS_st4_b9_c0 = nS_st3_b9_c0;
  assign nS_st4_b10_c0 = nS_st3_b10_c0;
  assign nS_st4_b11_c0 = nS_st3_b11_c0;
  assign nS_st4_b12_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b12_c0 : nS_st3_b12_c1;
  assign nS_st4_b13_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b13_c0 : nS_st3_b13_c1;
  assign nS_st4_b14_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b14_c0 : nS_st3_b14_c1;
  assign nS_st4_b15_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b15_c0 : nS_st3_b15_c1;
  assign nS_st4_b16_c0 = nS_st3_b16_c0;
  assign nS_st4_b17_c0 = nS_st3_b17_c0;
  assign nS_st4_b18_c0 = nS_st3_b18_c0;
  assign nS_st4_b19_c0 = nS_st3_b19_c0;
  assign nS_st4_b20_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b20_c0 : nS_st3_b20_c1;
  assign nS_st4_b21_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b21_c0 : nS_st3_b21_c1;
  assign nS_st4_b22_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b22_c0 : nS_st3_b22_c1;
  assign nS_st4_b23_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b23_c0 : nS_st3_b23_c1;
  assign nS_st4_b24_c0 = nS_st3_b24_c0;
  assign nS_st4_b25_c0 = nS_st3_b25_c0;
  assign nS_st4_b26_c0 = nS_st3_b26_c0;
  assign nS_st4_b27_c0 = nS_st3_b27_c0;
  assign nS_st4_b28_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b28_c0 : nS_st3_b28_c1;
  assign nS_st4_b29_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b29_c0 : nS_st3_b29_c1;
  assign nS_st4_b30_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b30_c0 : nS_st3_b30_c1;
  assign nS_st4_b31_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b31_c0 : nS_st3_b31_c1;
  assign nS_st4_b32_c0 = nS_st3_b32_c0;
  assign nS_st4_b33_c0 = nS_st3_b33_c0;
  assign nS_st4_b34_c0 = nS_st3_b34_c0;
  assign nS_st4_b35_c0 = nS_st3_b35_c0;
  assign nS_st4_b36_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b36_c0 : nS_st3_b36_c1;
  assign nS_st4_b37_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b37_c0 : nS_st3_b37_c1;
  assign nS_st4_b38_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b38_c0 : nS_st3_b38_c1;
  assign nS_st4_b39_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b39_c0 : nS_st3_b39_c1;
  assign nS_st4_b40_c0 = nS_st3_b40_c0;
  assign nS_st4_b41_c0 = nS_st3_b41_c0;
  assign nS_st4_b42_c0 = nS_st3_b42_c0;
  assign nS_st4_b43_c0 = nS_st3_b43_c0;
  assign nS_st4_b44_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b44_c0 : nS_st3_b44_c1;
  assign nS_st4_b45_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b45_c0 : nS_st3_b45_c1;
  assign nS_st4_b46_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b46_c0 : nS_st3_b46_c1;
  assign nS_st4_b47_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b47_c0 : nS_st3_b47_c1;
  assign nS_st4_b48_c0 = nS_st3_b48_c0;
  assign nS_st4_b49_c0 = nS_st3_b49_c0;
  assign nS_st4_b50_c0 = nS_st3_b50_c0;
  assign nS_st4_b51_c0 = nS_st3_b51_c0;
  assign nS_st4_b52_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b52_c0 : nS_st3_b52_c1;
  assign nS_st4_b53_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b53_c0 : nS_st3_b53_c1;
  assign nS_st4_b54_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b54_c0 : nS_st3_b54_c1;
  assign nS_st4_b55_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b55_c0 : nS_st3_b55_c1;
  assign nS_st4_b56_c0 = nS_st3_b56_c0;
  assign nS_st4_b57_c0 = nS_st3_b57_c0;
  assign nS_st4_b58_c0 = nS_st3_b58_c0;
  assign nS_st4_b59_c0 = nS_st3_b59_c0;
  assign nS_st4_b60_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b60_c0 : nS_st3_b60_c1;
  assign nS_st4_b61_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b61_c0 : nS_st3_b61_c1;
  assign nS_st4_b62_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b62_c0 : nS_st3_b62_c1;
  assign nS_st4_b63_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b63_c0 : nS_st3_b63_c1;
  assign nS_st4_b64_c0 = nS_st3_b64_c0;
  assign nS_st4_b65_c0 = nS_st3_b65_c0;
  assign nS_st4_b66_c0 = nS_st3_b66_c0;
  assign nS_st4_b67_c0 = nS_st3_b67_c0;
  assign nS_st4_b68_c0 = (nC_st3_b67_c0 == 0) ? nS_st3_b68_c0 : nS_st3_b68_c1;
  assign nS_st4_b69_c0 = (nC_st3_b67_c0 == 0) ? nS_st3_b69_c0 : nS_st3_b69_c1;
  assign nS_st4_b70_c0 = (nC_st3_b67_c0 == 0) ? nS_st3_b70_c0 : nS_st3_b70_c1;
  assign nS_st4_b71_c0 = (nC_st3_b67_c0 == 0) ? nS_st3_b71_c0 : nS_st3_b71_c1;
  assign nS_st4_b72_c0 = nS_st3_b72_c0;
  assign nS_st4_b73_c0 = nS_st3_b73_c0;
  assign nS_st4_b74_c0 = nS_st3_b74_c0;
  assign nS_st4_b75_c0 = nS_st3_b75_c0;
  assign nS_st4_b76_c0 = (nC_st3_b75_c0 == 0) ? nS_st3_b76_c0 : nS_st3_b76_c1;
  assign nS_st4_b77_c0 = (nC_st3_b75_c0 == 0) ? nS_st3_b77_c0 : nS_st3_b77_c1;
  assign nS_st4_b78_c0 = (nC_st3_b75_c0 == 0) ? nS_st3_b78_c0 : nS_st3_b78_c1;
  assign nS_st4_b79_c0 = (nC_st3_b75_c0 == 0) ? nS_st3_b79_c0 : nS_st3_b79_c1;
  assign nS_st4_b80_c0 = nS_st3_b80_c0;
  assign nS_st4_b81_c0 = nS_st3_b81_c0;
  assign nS_st4_b82_c0 = nS_st3_b82_c0;
  assign nS_st4_b83_c0 = nS_st3_b83_c0;
  assign nS_st4_b84_c0 = (nC_st3_b83_c0 == 0) ? nS_st3_b84_c0 : nS_st3_b84_c1;
  assign nS_st4_b85_c0 = (nC_st3_b83_c0 == 0) ? nS_st3_b85_c0 : nS_st3_b85_c1;
  assign nS_st4_b86_c0 = (nC_st3_b83_c0 == 0) ? nS_st3_b86_c0 : nS_st3_b86_c1;
  assign nS_st4_b87_c0 = (nC_st3_b83_c0 == 0) ? nS_st3_b87_c0 : nS_st3_b87_c1;
  assign nS_st4_b88_c0 = nS_st3_b88_c0;
  assign nS_st4_b89_c0 = nS_st3_b89_c0;
  assign nS_st4_b90_c0 = nS_st3_b90_c0;
  assign nS_st4_b91_c0 = nS_st3_b91_c0;
  assign nS_st4_b92_c0 = (nC_st3_b91_c0 == 0) ? nS_st3_b92_c0 : nS_st3_b92_c1;
  assign nS_st4_b93_c0 = (nC_st3_b91_c0 == 0) ? nS_st3_b93_c0 : nS_st3_b93_c1;
  assign nS_st4_b94_c0 = (nC_st3_b91_c0 == 0) ? nS_st3_b94_c0 : nS_st3_b94_c1;
  assign nS_st4_b95_c0 = (nC_st3_b91_c0 == 0) ? nS_st3_b95_c0 : nS_st3_b95_c1;
  assign nS_st4_b96_c0 = nS_st3_b96_c0;
  assign nS_st4_b97_c0 = nS_st3_b97_c0;
  assign nS_st4_b98_c0 = nS_st3_b98_c0;
  assign nS_st4_b99_c0 = nS_st3_b99_c0;
  assign nS_st4_b100_c0 = (nC_st3_b99_c0 == 0) ? nS_st3_b100_c0 : nS_st3_b100_c1;
  assign nS_st4_b101_c0 = (nC_st3_b99_c0 == 0) ? nS_st3_b101_c0 : nS_st3_b101_c1;
  assign nS_st4_b102_c0 = (nC_st3_b99_c0 == 0) ? nS_st3_b102_c0 : nS_st3_b102_c1;
  assign nS_st4_b103_c0 = (nC_st3_b99_c0 == 0) ? nS_st3_b103_c0 : nS_st3_b103_c1;
  assign nS_st4_b104_c0 = nS_st3_b104_c0;
  assign nS_st4_b105_c0 = nS_st3_b105_c0;
  assign nS_st4_b106_c0 = nS_st3_b106_c0;
  assign nS_st4_b107_c0 = nS_st3_b107_c0;
  assign nS_st4_b108_c0 = (nC_st3_b107_c0 == 0) ? nS_st3_b108_c0 : nS_st3_b108_c1;
  assign nS_st4_b109_c0 = (nC_st3_b107_c0 == 0) ? nS_st3_b109_c0 : nS_st3_b109_c1;
  assign nS_st4_b110_c0 = (nC_st3_b107_c0 == 0) ? nS_st3_b110_c0 : nS_st3_b110_c1;
  assign nS_st4_b111_c0 = (nC_st3_b107_c0 == 0) ? nS_st3_b111_c0 : nS_st3_b111_c1;
  assign nS_st4_b112_c0 = nS_st3_b112_c0;
  assign nS_st4_b113_c0 = nS_st3_b113_c0;
  assign nS_st4_b114_c0 = nS_st3_b114_c0;
  assign nS_st4_b115_c0 = nS_st3_b115_c0;
  assign nS_st4_b116_c0 = (nC_st3_b115_c0 == 0) ? nS_st3_b116_c0 : nS_st3_b116_c1;
  assign nS_st4_b117_c0 = (nC_st3_b115_c0 == 0) ? nS_st3_b117_c0 : nS_st3_b117_c1;
  assign nS_st4_b118_c0 = (nC_st3_b115_c0 == 0) ? nS_st3_b118_c0 : nS_st3_b118_c1;
  assign nS_st4_b119_c0 = (nC_st3_b115_c0 == 0) ? nS_st3_b119_c0 : nS_st3_b119_c1;
  assign nS_st4_b120_c0 = nS_st3_b120_c0;
  assign nS_st4_b121_c0 = nS_st3_b121_c0;
  assign nS_st4_b122_c0 = nS_st3_b122_c0;
  assign nS_st4_b123_c0 = nS_st3_b123_c0;
  assign nS_st4_b124_c0 = (nC_st3_b123_c0 == 0) ? nS_st3_b124_c0 : nS_st3_b124_c1;
  assign nS_st4_b125_c0 = (nC_st3_b123_c0 == 0) ? nS_st3_b125_c0 : nS_st3_b125_c1;
  assign nS_st4_b126_c0 = (nC_st3_b123_c0 == 0) ? nS_st3_b126_c0 : nS_st3_b126_c1;
  assign nS_st4_b127_c0 = (nC_st3_b123_c0 == 0) ? nS_st3_b127_c0 : nS_st3_b127_c1;
  assign nS_st4_b0_c1 = nS_st3_b0_c1;
  assign nS_st4_b1_c1 = nS_st3_b1_c1;
  assign nS_st4_b2_c1 = nS_st3_b2_c1;
  assign nS_st4_b3_c1 = nS_st3_b3_c1;
  assign nS_st4_b4_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b4_c0 : nS_st3_b4_c1;
  assign nS_st4_b5_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b5_c0 : nS_st3_b5_c1;
  assign nS_st4_b6_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b6_c0 : nS_st3_b6_c1;
  assign nS_st4_b7_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b7_c0 : nS_st3_b7_c1;
  assign nS_st4_b8_c1 = nS_st3_b8_c1;
  assign nS_st4_b9_c1 = nS_st3_b9_c1;
  assign nS_st4_b10_c1 = nS_st3_b10_c1;
  assign nS_st4_b11_c1 = nS_st3_b11_c1;
  assign nS_st4_b12_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b12_c0 : nS_st3_b12_c1;
  assign nS_st4_b13_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b13_c0 : nS_st3_b13_c1;
  assign nS_st4_b14_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b14_c0 : nS_st3_b14_c1;
  assign nS_st4_b15_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b15_c0 : nS_st3_b15_c1;
  assign nS_st4_b16_c1 = nS_st3_b16_c1;
  assign nS_st4_b17_c1 = nS_st3_b17_c1;
  assign nS_st4_b18_c1 = nS_st3_b18_c1;
  assign nS_st4_b19_c1 = nS_st3_b19_c1;
  assign nS_st4_b20_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b20_c0 : nS_st3_b20_c1;
  assign nS_st4_b21_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b21_c0 : nS_st3_b21_c1;
  assign nS_st4_b22_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b22_c0 : nS_st3_b22_c1;
  assign nS_st4_b23_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b23_c0 : nS_st3_b23_c1;
  assign nS_st4_b24_c1 = nS_st3_b24_c1;
  assign nS_st4_b25_c1 = nS_st3_b25_c1;
  assign nS_st4_b26_c1 = nS_st3_b26_c1;
  assign nS_st4_b27_c1 = nS_st3_b27_c1;
  assign nS_st4_b28_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b28_c0 : nS_st3_b28_c1;
  assign nS_st4_b29_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b29_c0 : nS_st3_b29_c1;
  assign nS_st4_b30_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b30_c0 : nS_st3_b30_c1;
  assign nS_st4_b31_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b31_c0 : nS_st3_b31_c1;
  assign nS_st4_b32_c1 = nS_st3_b32_c1;
  assign nS_st4_b33_c1 = nS_st3_b33_c1;
  assign nS_st4_b34_c1 = nS_st3_b34_c1;
  assign nS_st4_b35_c1 = nS_st3_b35_c1;
  assign nS_st4_b36_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b36_c0 : nS_st3_b36_c1;
  assign nS_st4_b37_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b37_c0 : nS_st3_b37_c1;
  assign nS_st4_b38_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b38_c0 : nS_st3_b38_c1;
  assign nS_st4_b39_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b39_c0 : nS_st3_b39_c1;
  assign nS_st4_b40_c1 = nS_st3_b40_c1;
  assign nS_st4_b41_c1 = nS_st3_b41_c1;
  assign nS_st4_b42_c1 = nS_st3_b42_c1;
  assign nS_st4_b43_c1 = nS_st3_b43_c1;
  assign nS_st4_b44_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b44_c0 : nS_st3_b44_c1;
  assign nS_st4_b45_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b45_c0 : nS_st3_b45_c1;
  assign nS_st4_b46_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b46_c0 : nS_st3_b46_c1;
  assign nS_st4_b47_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b47_c0 : nS_st3_b47_c1;
  assign nS_st4_b48_c1 = nS_st3_b48_c1;
  assign nS_st4_b49_c1 = nS_st3_b49_c1;
  assign nS_st4_b50_c1 = nS_st3_b50_c1;
  assign nS_st4_b51_c1 = nS_st3_b51_c1;
  assign nS_st4_b52_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b52_c0 : nS_st3_b52_c1;
  assign nS_st4_b53_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b53_c0 : nS_st3_b53_c1;
  assign nS_st4_b54_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b54_c0 : nS_st3_b54_c1;
  assign nS_st4_b55_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b55_c0 : nS_st3_b55_c1;
  assign nS_st4_b56_c1 = nS_st3_b56_c1;
  assign nS_st4_b57_c1 = nS_st3_b57_c1;
  assign nS_st4_b58_c1 = nS_st3_b58_c1;
  assign nS_st4_b59_c1 = nS_st3_b59_c1;
  assign nS_st4_b60_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b60_c0 : nS_st3_b60_c1;
  assign nS_st4_b61_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b61_c0 : nS_st3_b61_c1;
  assign nS_st4_b62_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b62_c0 : nS_st3_b62_c1;
  assign nS_st4_b63_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b63_c0 : nS_st3_b63_c1;
  assign nS_st4_b64_c1 = nS_st3_b64_c1;
  assign nS_st4_b65_c1 = nS_st3_b65_c1;
  assign nS_st4_b66_c1 = nS_st3_b66_c1;
  assign nS_st4_b67_c1 = nS_st3_b67_c1;
  assign nS_st4_b68_c1 = (nC_st3_b67_c1 == 0) ? nS_st3_b68_c0 : nS_st3_b68_c1;
  assign nS_st4_b69_c1 = (nC_st3_b67_c1 == 0) ? nS_st3_b69_c0 : nS_st3_b69_c1;
  assign nS_st4_b70_c1 = (nC_st3_b67_c1 == 0) ? nS_st3_b70_c0 : nS_st3_b70_c1;
  assign nS_st4_b71_c1 = (nC_st3_b67_c1 == 0) ? nS_st3_b71_c0 : nS_st3_b71_c1;
  assign nS_st4_b72_c1 = nS_st3_b72_c1;
  assign nS_st4_b73_c1 = nS_st3_b73_c1;
  assign nS_st4_b74_c1 = nS_st3_b74_c1;
  assign nS_st4_b75_c1 = nS_st3_b75_c1;
  assign nS_st4_b76_c1 = (nC_st3_b75_c1 == 0) ? nS_st3_b76_c0 : nS_st3_b76_c1;
  assign nS_st4_b77_c1 = (nC_st3_b75_c1 == 0) ? nS_st3_b77_c0 : nS_st3_b77_c1;
  assign nS_st4_b78_c1 = (nC_st3_b75_c1 == 0) ? nS_st3_b78_c0 : nS_st3_b78_c1;
  assign nS_st4_b79_c1 = (nC_st3_b75_c1 == 0) ? nS_st3_b79_c0 : nS_st3_b79_c1;
  assign nS_st4_b80_c1 = nS_st3_b80_c1;
  assign nS_st4_b81_c1 = nS_st3_b81_c1;
  assign nS_st4_b82_c1 = nS_st3_b82_c1;
  assign nS_st4_b83_c1 = nS_st3_b83_c1;
  assign nS_st4_b84_c1 = (nC_st3_b83_c1 == 0) ? nS_st3_b84_c0 : nS_st3_b84_c1;
  assign nS_st4_b85_c1 = (nC_st3_b83_c1 == 0) ? nS_st3_b85_c0 : nS_st3_b85_c1;
  assign nS_st4_b86_c1 = (nC_st3_b83_c1 == 0) ? nS_st3_b86_c0 : nS_st3_b86_c1;
  assign nS_st4_b87_c1 = (nC_st3_b83_c1 == 0) ? nS_st3_b87_c0 : nS_st3_b87_c1;
  assign nS_st4_b88_c1 = nS_st3_b88_c1;
  assign nS_st4_b89_c1 = nS_st3_b89_c1;
  assign nS_st4_b90_c1 = nS_st3_b90_c1;
  assign nS_st4_b91_c1 = nS_st3_b91_c1;
  assign nS_st4_b92_c1 = (nC_st3_b91_c1 == 0) ? nS_st3_b92_c0 : nS_st3_b92_c1;
  assign nS_st4_b93_c1 = (nC_st3_b91_c1 == 0) ? nS_st3_b93_c0 : nS_st3_b93_c1;
  assign nS_st4_b94_c1 = (nC_st3_b91_c1 == 0) ? nS_st3_b94_c0 : nS_st3_b94_c1;
  assign nS_st4_b95_c1 = (nC_st3_b91_c1 == 0) ? nS_st3_b95_c0 : nS_st3_b95_c1;
  assign nS_st4_b96_c1 = nS_st3_b96_c1;
  assign nS_st4_b97_c1 = nS_st3_b97_c1;
  assign nS_st4_b98_c1 = nS_st3_b98_c1;
  assign nS_st4_b99_c1 = nS_st3_b99_c1;
  assign nS_st4_b100_c1 = (nC_st3_b99_c1 == 0) ? nS_st3_b100_c0 : nS_st3_b100_c1;
  assign nS_st4_b101_c1 = (nC_st3_b99_c1 == 0) ? nS_st3_b101_c0 : nS_st3_b101_c1;
  assign nS_st4_b102_c1 = (nC_st3_b99_c1 == 0) ? nS_st3_b102_c0 : nS_st3_b102_c1;
  assign nS_st4_b103_c1 = (nC_st3_b99_c1 == 0) ? nS_st3_b103_c0 : nS_st3_b103_c1;
  assign nS_st4_b104_c1 = nS_st3_b104_c1;
  assign nS_st4_b105_c1 = nS_st3_b105_c1;
  assign nS_st4_b106_c1 = nS_st3_b106_c1;
  assign nS_st4_b107_c1 = nS_st3_b107_c1;
  assign nS_st4_b108_c1 = (nC_st3_b107_c1 == 0) ? nS_st3_b108_c0 : nS_st3_b108_c1;
  assign nS_st4_b109_c1 = (nC_st3_b107_c1 == 0) ? nS_st3_b109_c0 : nS_st3_b109_c1;
  assign nS_st4_b110_c1 = (nC_st3_b107_c1 == 0) ? nS_st3_b110_c0 : nS_st3_b110_c1;
  assign nS_st4_b111_c1 = (nC_st3_b107_c1 == 0) ? nS_st3_b111_c0 : nS_st3_b111_c1;
  assign nS_st4_b112_c1 = nS_st3_b112_c1;
  assign nS_st4_b113_c1 = nS_st3_b113_c1;
  assign nS_st4_b114_c1 = nS_st3_b114_c1;
  assign nS_st4_b115_c1 = nS_st3_b115_c1;
  assign nS_st4_b116_c1 = (nC_st3_b115_c1 == 0) ? nS_st3_b116_c0 : nS_st3_b116_c1;
  assign nS_st4_b117_c1 = (nC_st3_b115_c1 == 0) ? nS_st3_b117_c0 : nS_st3_b117_c1;
  assign nS_st4_b118_c1 = (nC_st3_b115_c1 == 0) ? nS_st3_b118_c0 : nS_st3_b118_c1;
  assign nS_st4_b119_c1 = (nC_st3_b115_c1 == 0) ? nS_st3_b119_c0 : nS_st3_b119_c1;
  assign nS_st4_b120_c1 = nS_st3_b120_c1;
  assign nS_st4_b121_c1 = nS_st3_b121_c1;
  assign nS_st4_b122_c1 = nS_st3_b122_c1;
  assign nS_st4_b123_c1 = nS_st3_b123_c1;
  assign nS_st4_b124_c1 = (nC_st3_b123_c1 == 0) ? nS_st3_b124_c0 : nS_st3_b124_c1;
  assign nS_st4_b125_c1 = (nC_st3_b123_c1 == 0) ? nS_st3_b125_c0 : nS_st3_b125_c1;
  assign nS_st4_b126_c1 = (nC_st3_b123_c1 == 0) ? nS_st3_b126_c0 : nS_st3_b126_c1;
  assign nS_st4_b127_c1 = (nC_st3_b123_c1 == 0) ? nS_st3_b127_c0 : nS_st3_b127_c1;
  assign nC_st4_b7_c0 = (nC_st3_b3_c0 == 0) ? nC_st3_b7_c0 : nC_st3_b7_c1;
  assign nC_st4_b15_c0 = (nC_st3_b11_c0 == 0) ? nC_st3_b15_c0 : nC_st3_b15_c1;
  assign nC_st4_b23_c0 = (nC_st3_b19_c0 == 0) ? nC_st3_b23_c0 : nC_st3_b23_c1;
  assign nC_st4_b31_c0 = (nC_st3_b27_c0 == 0) ? nC_st3_b31_c0 : nC_st3_b31_c1;
  assign nC_st4_b39_c0 = (nC_st3_b35_c0 == 0) ? nC_st3_b39_c0 : nC_st3_b39_c1;
  assign nC_st4_b47_c0 = (nC_st3_b43_c0 == 0) ? nC_st3_b47_c0 : nC_st3_b47_c1;
  assign nC_st4_b55_c0 = (nC_st3_b51_c0 == 0) ? nC_st3_b55_c0 : nC_st3_b55_c1;
  assign nC_st4_b63_c0 = (nC_st3_b59_c0 == 0) ? nC_st3_b63_c0 : nC_st3_b63_c1;
  assign nC_st4_b71_c0 = (nC_st3_b67_c0 == 0) ? nC_st3_b71_c0 : nC_st3_b71_c1;
  assign nC_st4_b79_c0 = (nC_st3_b75_c0 == 0) ? nC_st3_b79_c0 : nC_st3_b79_c1;
  assign nC_st4_b87_c0 = (nC_st3_b83_c0 == 0) ? nC_st3_b87_c0 : nC_st3_b87_c1;
  assign nC_st4_b95_c0 = (nC_st3_b91_c0 == 0) ? nC_st3_b95_c0 : nC_st3_b95_c1;
  assign nC_st4_b103_c0 = (nC_st3_b99_c0 == 0) ? nC_st3_b103_c0 : nC_st3_b103_c1;
  assign nC_st4_b111_c0 = (nC_st3_b107_c0 == 0) ? nC_st3_b111_c0 : nC_st3_b111_c1;
  assign nC_st4_b119_c0 = (nC_st3_b115_c0 == 0) ? nC_st3_b119_c0 : nC_st3_b119_c1;
  assign nC_st4_b127_c0 = (nC_st3_b123_c0 == 0) ? nC_st3_b127_c0 : nC_st3_b127_c1;
  assign nC_st4_b7_c1 = (nC_st3_b3_c1 == 0) ? nC_st3_b7_c0 : nC_st3_b7_c1;
  assign nC_st4_b15_c1 = (nC_st3_b11_c1 == 0) ? nC_st3_b15_c0 : nC_st3_b15_c1;
  assign nC_st4_b23_c1 = (nC_st3_b19_c1 == 0) ? nC_st3_b23_c0 : nC_st3_b23_c1;
  assign nC_st4_b31_c1 = (nC_st3_b27_c1 == 0) ? nC_st3_b31_c0 : nC_st3_b31_c1;
  assign nC_st4_b39_c1 = (nC_st3_b35_c1 == 0) ? nC_st3_b39_c0 : nC_st3_b39_c1;
  assign nC_st4_b47_c1 = (nC_st3_b43_c1 == 0) ? nC_st3_b47_c0 : nC_st3_b47_c1;
  assign nC_st4_b55_c1 = (nC_st3_b51_c1 == 0) ? nC_st3_b55_c0 : nC_st3_b55_c1;
  assign nC_st4_b63_c1 = (nC_st3_b59_c1 == 0) ? nC_st3_b63_c0 : nC_st3_b63_c1;
  assign nC_st4_b71_c1 = (nC_st3_b67_c1 == 0) ? nC_st3_b71_c0 : nC_st3_b71_c1;
  assign nC_st4_b79_c1 = (nC_st3_b75_c1 == 0) ? nC_st3_b79_c0 : nC_st3_b79_c1;
  assign nC_st4_b87_c1 = (nC_st3_b83_c1 == 0) ? nC_st3_b87_c0 : nC_st3_b87_c1;
  assign nC_st4_b95_c1 = (nC_st3_b91_c1 == 0) ? nC_st3_b95_c0 : nC_st3_b95_c1;
  assign nC_st4_b103_c1 = (nC_st3_b99_c1 == 0) ? nC_st3_b103_c0 : nC_st3_b103_c1;
  assign nC_st4_b111_c1 = (nC_st3_b107_c1 == 0) ? nC_st3_b111_c0 : nC_st3_b111_c1;
  assign nC_st4_b119_c1 = (nC_st3_b115_c1 == 0) ? nC_st3_b119_c0 : nC_st3_b119_c1;
  assign nC_st4_b127_c1 = (nC_st3_b123_c1 == 0) ? nC_st3_b127_c0 : nC_st3_b127_c1;

  assign nS_st5_b0_c0 = nS_st4_b0_c0;
  assign nS_st5_b1_c0 = nS_st4_b1_c0;
  assign nS_st5_b2_c0 = nS_st4_b2_c0;
  assign nS_st5_b3_c0 = nS_st4_b3_c0;
  assign nS_st5_b4_c0 = nS_st4_b4_c0;
  assign nS_st5_b5_c0 = nS_st4_b5_c0;
  assign nS_st5_b6_c0 = nS_st4_b6_c0;
  assign nS_st5_b7_c0 = nS_st4_b7_c0;
  assign nS_st5_b8_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b8_c0 : nS_st4_b8_c1;
  assign nS_st5_b9_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b9_c0 : nS_st4_b9_c1;
  assign nS_st5_b10_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b10_c0 : nS_st4_b10_c1;
  assign nS_st5_b11_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b11_c0 : nS_st4_b11_c1;
  assign nS_st5_b12_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b12_c0 : nS_st4_b12_c1;
  assign nS_st5_b13_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b13_c0 : nS_st4_b13_c1;
  assign nS_st5_b14_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b14_c0 : nS_st4_b14_c1;
  assign nS_st5_b15_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b15_c0 : nS_st4_b15_c1;
  assign nS_st5_b16_c0 = nS_st4_b16_c0;
  assign nS_st5_b17_c0 = nS_st4_b17_c0;
  assign nS_st5_b18_c0 = nS_st4_b18_c0;
  assign nS_st5_b19_c0 = nS_st4_b19_c0;
  assign nS_st5_b20_c0 = nS_st4_b20_c0;
  assign nS_st5_b21_c0 = nS_st4_b21_c0;
  assign nS_st5_b22_c0 = nS_st4_b22_c0;
  assign nS_st5_b23_c0 = nS_st4_b23_c0;
  assign nS_st5_b24_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b24_c0 : nS_st4_b24_c1;
  assign nS_st5_b25_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b25_c0 : nS_st4_b25_c1;
  assign nS_st5_b26_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b26_c0 : nS_st4_b26_c1;
  assign nS_st5_b27_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b27_c0 : nS_st4_b27_c1;
  assign nS_st5_b28_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b28_c0 : nS_st4_b28_c1;
  assign nS_st5_b29_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b29_c0 : nS_st4_b29_c1;
  assign nS_st5_b30_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b30_c0 : nS_st4_b30_c1;
  assign nS_st5_b31_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b31_c0 : nS_st4_b31_c1;
  assign nS_st5_b32_c0 = nS_st4_b32_c0;
  assign nS_st5_b33_c0 = nS_st4_b33_c0;
  assign nS_st5_b34_c0 = nS_st4_b34_c0;
  assign nS_st5_b35_c0 = nS_st4_b35_c0;
  assign nS_st5_b36_c0 = nS_st4_b36_c0;
  assign nS_st5_b37_c0 = nS_st4_b37_c0;
  assign nS_st5_b38_c0 = nS_st4_b38_c0;
  assign nS_st5_b39_c0 = nS_st4_b39_c0;
  assign nS_st5_b40_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b40_c0 : nS_st4_b40_c1;
  assign nS_st5_b41_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b41_c0 : nS_st4_b41_c1;
  assign nS_st5_b42_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b42_c0 : nS_st4_b42_c1;
  assign nS_st5_b43_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b43_c0 : nS_st4_b43_c1;
  assign nS_st5_b44_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b44_c0 : nS_st4_b44_c1;
  assign nS_st5_b45_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b45_c0 : nS_st4_b45_c1;
  assign nS_st5_b46_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b46_c0 : nS_st4_b46_c1;
  assign nS_st5_b47_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b47_c0 : nS_st4_b47_c1;
  assign nS_st5_b48_c0 = nS_st4_b48_c0;
  assign nS_st5_b49_c0 = nS_st4_b49_c0;
  assign nS_st5_b50_c0 = nS_st4_b50_c0;
  assign nS_st5_b51_c0 = nS_st4_b51_c0;
  assign nS_st5_b52_c0 = nS_st4_b52_c0;
  assign nS_st5_b53_c0 = nS_st4_b53_c0;
  assign nS_st5_b54_c0 = nS_st4_b54_c0;
  assign nS_st5_b55_c0 = nS_st4_b55_c0;
  assign nS_st5_b56_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b56_c0 : nS_st4_b56_c1;
  assign nS_st5_b57_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b57_c0 : nS_st4_b57_c1;
  assign nS_st5_b58_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b58_c0 : nS_st4_b58_c1;
  assign nS_st5_b59_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b59_c0 : nS_st4_b59_c1;
  assign nS_st5_b60_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b60_c0 : nS_st4_b60_c1;
  assign nS_st5_b61_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b61_c0 : nS_st4_b61_c1;
  assign nS_st5_b62_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b62_c0 : nS_st4_b62_c1;
  assign nS_st5_b63_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b63_c0 : nS_st4_b63_c1;
  assign nS_st5_b64_c0 = nS_st4_b64_c0;
  assign nS_st5_b65_c0 = nS_st4_b65_c0;
  assign nS_st5_b66_c0 = nS_st4_b66_c0;
  assign nS_st5_b67_c0 = nS_st4_b67_c0;
  assign nS_st5_b68_c0 = nS_st4_b68_c0;
  assign nS_st5_b69_c0 = nS_st4_b69_c0;
  assign nS_st5_b70_c0 = nS_st4_b70_c0;
  assign nS_st5_b71_c0 = nS_st4_b71_c0;
  assign nS_st5_b72_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b72_c0 : nS_st4_b72_c1;
  assign nS_st5_b73_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b73_c0 : nS_st4_b73_c1;
  assign nS_st5_b74_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b74_c0 : nS_st4_b74_c1;
  assign nS_st5_b75_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b75_c0 : nS_st4_b75_c1;
  assign nS_st5_b76_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b76_c0 : nS_st4_b76_c1;
  assign nS_st5_b77_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b77_c0 : nS_st4_b77_c1;
  assign nS_st5_b78_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b78_c0 : nS_st4_b78_c1;
  assign nS_st5_b79_c0 = (nC_st4_b71_c0 == 0) ? nS_st4_b79_c0 : nS_st4_b79_c1;
  assign nS_st5_b80_c0 = nS_st4_b80_c0;
  assign nS_st5_b81_c0 = nS_st4_b81_c0;
  assign nS_st5_b82_c0 = nS_st4_b82_c0;
  assign nS_st5_b83_c0 = nS_st4_b83_c0;
  assign nS_st5_b84_c0 = nS_st4_b84_c0;
  assign nS_st5_b85_c0 = nS_st4_b85_c0;
  assign nS_st5_b86_c0 = nS_st4_b86_c0;
  assign nS_st5_b87_c0 = nS_st4_b87_c0;
  assign nS_st5_b88_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b88_c0 : nS_st4_b88_c1;
  assign nS_st5_b89_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b89_c0 : nS_st4_b89_c1;
  assign nS_st5_b90_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b90_c0 : nS_st4_b90_c1;
  assign nS_st5_b91_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b91_c0 : nS_st4_b91_c1;
  assign nS_st5_b92_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b92_c0 : nS_st4_b92_c1;
  assign nS_st5_b93_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b93_c0 : nS_st4_b93_c1;
  assign nS_st5_b94_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b94_c0 : nS_st4_b94_c1;
  assign nS_st5_b95_c0 = (nC_st4_b87_c0 == 0) ? nS_st4_b95_c0 : nS_st4_b95_c1;
  assign nS_st5_b96_c0 = nS_st4_b96_c0;
  assign nS_st5_b97_c0 = nS_st4_b97_c0;
  assign nS_st5_b98_c0 = nS_st4_b98_c0;
  assign nS_st5_b99_c0 = nS_st4_b99_c0;
  assign nS_st5_b100_c0 = nS_st4_b100_c0;
  assign nS_st5_b101_c0 = nS_st4_b101_c0;
  assign nS_st5_b102_c0 = nS_st4_b102_c0;
  assign nS_st5_b103_c0 = nS_st4_b103_c0;
  assign nS_st5_b104_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b104_c0 : nS_st4_b104_c1;
  assign nS_st5_b105_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b105_c0 : nS_st4_b105_c1;
  assign nS_st5_b106_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b106_c0 : nS_st4_b106_c1;
  assign nS_st5_b107_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b107_c0 : nS_st4_b107_c1;
  assign nS_st5_b108_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b108_c0 : nS_st4_b108_c1;
  assign nS_st5_b109_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b109_c0 : nS_st4_b109_c1;
  assign nS_st5_b110_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b110_c0 : nS_st4_b110_c1;
  assign nS_st5_b111_c0 = (nC_st4_b103_c0 == 0) ? nS_st4_b111_c0 : nS_st4_b111_c1;
  assign nS_st5_b112_c0 = nS_st4_b112_c0;
  assign nS_st5_b113_c0 = nS_st4_b113_c0;
  assign nS_st5_b114_c0 = nS_st4_b114_c0;
  assign nS_st5_b115_c0 = nS_st4_b115_c0;
  assign nS_st5_b116_c0 = nS_st4_b116_c0;
  assign nS_st5_b117_c0 = nS_st4_b117_c0;
  assign nS_st5_b118_c0 = nS_st4_b118_c0;
  assign nS_st5_b119_c0 = nS_st4_b119_c0;
  assign nS_st5_b120_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b120_c0 : nS_st4_b120_c1;
  assign nS_st5_b121_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b121_c0 : nS_st4_b121_c1;
  assign nS_st5_b122_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b122_c0 : nS_st4_b122_c1;
  assign nS_st5_b123_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b123_c0 : nS_st4_b123_c1;
  assign nS_st5_b124_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b124_c0 : nS_st4_b124_c1;
  assign nS_st5_b125_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b125_c0 : nS_st4_b125_c1;
  assign nS_st5_b126_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b126_c0 : nS_st4_b126_c1;
  assign nS_st5_b127_c0 = (nC_st4_b119_c0 == 0) ? nS_st4_b127_c0 : nS_st4_b127_c1;
  assign nS_st5_b0_c1 = nS_st4_b0_c1;
  assign nS_st5_b1_c1 = nS_st4_b1_c1;
  assign nS_st5_b2_c1 = nS_st4_b2_c1;
  assign nS_st5_b3_c1 = nS_st4_b3_c1;
  assign nS_st5_b4_c1 = nS_st4_b4_c1;
  assign nS_st5_b5_c1 = nS_st4_b5_c1;
  assign nS_st5_b6_c1 = nS_st4_b6_c1;
  assign nS_st5_b7_c1 = nS_st4_b7_c1;
  assign nS_st5_b8_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b8_c0 : nS_st4_b8_c1;
  assign nS_st5_b9_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b9_c0 : nS_st4_b9_c1;
  assign nS_st5_b10_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b10_c0 : nS_st4_b10_c1;
  assign nS_st5_b11_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b11_c0 : nS_st4_b11_c1;
  assign nS_st5_b12_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b12_c0 : nS_st4_b12_c1;
  assign nS_st5_b13_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b13_c0 : nS_st4_b13_c1;
  assign nS_st5_b14_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b14_c0 : nS_st4_b14_c1;
  assign nS_st5_b15_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b15_c0 : nS_st4_b15_c1;
  assign nS_st5_b16_c1 = nS_st4_b16_c1;
  assign nS_st5_b17_c1 = nS_st4_b17_c1;
  assign nS_st5_b18_c1 = nS_st4_b18_c1;
  assign nS_st5_b19_c1 = nS_st4_b19_c1;
  assign nS_st5_b20_c1 = nS_st4_b20_c1;
  assign nS_st5_b21_c1 = nS_st4_b21_c1;
  assign nS_st5_b22_c1 = nS_st4_b22_c1;
  assign nS_st5_b23_c1 = nS_st4_b23_c1;
  assign nS_st5_b24_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b24_c0 : nS_st4_b24_c1;
  assign nS_st5_b25_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b25_c0 : nS_st4_b25_c1;
  assign nS_st5_b26_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b26_c0 : nS_st4_b26_c1;
  assign nS_st5_b27_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b27_c0 : nS_st4_b27_c1;
  assign nS_st5_b28_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b28_c0 : nS_st4_b28_c1;
  assign nS_st5_b29_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b29_c0 : nS_st4_b29_c1;
  assign nS_st5_b30_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b30_c0 : nS_st4_b30_c1;
  assign nS_st5_b31_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b31_c0 : nS_st4_b31_c1;
  assign nS_st5_b32_c1 = nS_st4_b32_c1;
  assign nS_st5_b33_c1 = nS_st4_b33_c1;
  assign nS_st5_b34_c1 = nS_st4_b34_c1;
  assign nS_st5_b35_c1 = nS_st4_b35_c1;
  assign nS_st5_b36_c1 = nS_st4_b36_c1;
  assign nS_st5_b37_c1 = nS_st4_b37_c1;
  assign nS_st5_b38_c1 = nS_st4_b38_c1;
  assign nS_st5_b39_c1 = nS_st4_b39_c1;
  assign nS_st5_b40_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b40_c0 : nS_st4_b40_c1;
  assign nS_st5_b41_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b41_c0 : nS_st4_b41_c1;
  assign nS_st5_b42_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b42_c0 : nS_st4_b42_c1;
  assign nS_st5_b43_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b43_c0 : nS_st4_b43_c1;
  assign nS_st5_b44_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b44_c0 : nS_st4_b44_c1;
  assign nS_st5_b45_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b45_c0 : nS_st4_b45_c1;
  assign nS_st5_b46_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b46_c0 : nS_st4_b46_c1;
  assign nS_st5_b47_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b47_c0 : nS_st4_b47_c1;
  assign nS_st5_b48_c1 = nS_st4_b48_c1;
  assign nS_st5_b49_c1 = nS_st4_b49_c1;
  assign nS_st5_b50_c1 = nS_st4_b50_c1;
  assign nS_st5_b51_c1 = nS_st4_b51_c1;
  assign nS_st5_b52_c1 = nS_st4_b52_c1;
  assign nS_st5_b53_c1 = nS_st4_b53_c1;
  assign nS_st5_b54_c1 = nS_st4_b54_c1;
  assign nS_st5_b55_c1 = nS_st4_b55_c1;
  assign nS_st5_b56_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b56_c0 : nS_st4_b56_c1;
  assign nS_st5_b57_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b57_c0 : nS_st4_b57_c1;
  assign nS_st5_b58_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b58_c0 : nS_st4_b58_c1;
  assign nS_st5_b59_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b59_c0 : nS_st4_b59_c1;
  assign nS_st5_b60_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b60_c0 : nS_st4_b60_c1;
  assign nS_st5_b61_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b61_c0 : nS_st4_b61_c1;
  assign nS_st5_b62_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b62_c0 : nS_st4_b62_c1;
  assign nS_st5_b63_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b63_c0 : nS_st4_b63_c1;
  assign nS_st5_b64_c1 = nS_st4_b64_c1;
  assign nS_st5_b65_c1 = nS_st4_b65_c1;
  assign nS_st5_b66_c1 = nS_st4_b66_c1;
  assign nS_st5_b67_c1 = nS_st4_b67_c1;
  assign nS_st5_b68_c1 = nS_st4_b68_c1;
  assign nS_st5_b69_c1 = nS_st4_b69_c1;
  assign nS_st5_b70_c1 = nS_st4_b70_c1;
  assign nS_st5_b71_c1 = nS_st4_b71_c1;
  assign nS_st5_b72_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b72_c0 : nS_st4_b72_c1;
  assign nS_st5_b73_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b73_c0 : nS_st4_b73_c1;
  assign nS_st5_b74_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b74_c0 : nS_st4_b74_c1;
  assign nS_st5_b75_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b75_c0 : nS_st4_b75_c1;
  assign nS_st5_b76_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b76_c0 : nS_st4_b76_c1;
  assign nS_st5_b77_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b77_c0 : nS_st4_b77_c1;
  assign nS_st5_b78_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b78_c0 : nS_st4_b78_c1;
  assign nS_st5_b79_c1 = (nC_st4_b71_c1 == 0) ? nS_st4_b79_c0 : nS_st4_b79_c1;
  assign nS_st5_b80_c1 = nS_st4_b80_c1;
  assign nS_st5_b81_c1 = nS_st4_b81_c1;
  assign nS_st5_b82_c1 = nS_st4_b82_c1;
  assign nS_st5_b83_c1 = nS_st4_b83_c1;
  assign nS_st5_b84_c1 = nS_st4_b84_c1;
  assign nS_st5_b85_c1 = nS_st4_b85_c1;
  assign nS_st5_b86_c1 = nS_st4_b86_c1;
  assign nS_st5_b87_c1 = nS_st4_b87_c1;
  assign nS_st5_b88_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b88_c0 : nS_st4_b88_c1;
  assign nS_st5_b89_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b89_c0 : nS_st4_b89_c1;
  assign nS_st5_b90_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b90_c0 : nS_st4_b90_c1;
  assign nS_st5_b91_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b91_c0 : nS_st4_b91_c1;
  assign nS_st5_b92_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b92_c0 : nS_st4_b92_c1;
  assign nS_st5_b93_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b93_c0 : nS_st4_b93_c1;
  assign nS_st5_b94_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b94_c0 : nS_st4_b94_c1;
  assign nS_st5_b95_c1 = (nC_st4_b87_c1 == 0) ? nS_st4_b95_c0 : nS_st4_b95_c1;
  assign nS_st5_b96_c1 = nS_st4_b96_c1;
  assign nS_st5_b97_c1 = nS_st4_b97_c1;
  assign nS_st5_b98_c1 = nS_st4_b98_c1;
  assign nS_st5_b99_c1 = nS_st4_b99_c1;
  assign nS_st5_b100_c1 = nS_st4_b100_c1;
  assign nS_st5_b101_c1 = nS_st4_b101_c1;
  assign nS_st5_b102_c1 = nS_st4_b102_c1;
  assign nS_st5_b103_c1 = nS_st4_b103_c1;
  assign nS_st5_b104_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b104_c0 : nS_st4_b104_c1;
  assign nS_st5_b105_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b105_c0 : nS_st4_b105_c1;
  assign nS_st5_b106_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b106_c0 : nS_st4_b106_c1;
  assign nS_st5_b107_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b107_c0 : nS_st4_b107_c1;
  assign nS_st5_b108_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b108_c0 : nS_st4_b108_c1;
  assign nS_st5_b109_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b109_c0 : nS_st4_b109_c1;
  assign nS_st5_b110_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b110_c0 : nS_st4_b110_c1;
  assign nS_st5_b111_c1 = (nC_st4_b103_c1 == 0) ? nS_st4_b111_c0 : nS_st4_b111_c1;
  assign nS_st5_b112_c1 = nS_st4_b112_c1;
  assign nS_st5_b113_c1 = nS_st4_b113_c1;
  assign nS_st5_b114_c1 = nS_st4_b114_c1;
  assign nS_st5_b115_c1 = nS_st4_b115_c1;
  assign nS_st5_b116_c1 = nS_st4_b116_c1;
  assign nS_st5_b117_c1 = nS_st4_b117_c1;
  assign nS_st5_b118_c1 = nS_st4_b118_c1;
  assign nS_st5_b119_c1 = nS_st4_b119_c1;
  assign nS_st5_b120_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b120_c0 : nS_st4_b120_c1;
  assign nS_st5_b121_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b121_c0 : nS_st4_b121_c1;
  assign nS_st5_b122_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b122_c0 : nS_st4_b122_c1;
  assign nS_st5_b123_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b123_c0 : nS_st4_b123_c1;
  assign nS_st5_b124_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b124_c0 : nS_st4_b124_c1;
  assign nS_st5_b125_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b125_c0 : nS_st4_b125_c1;
  assign nS_st5_b126_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b126_c0 : nS_st4_b126_c1;
  assign nS_st5_b127_c1 = (nC_st4_b119_c1 == 0) ? nS_st4_b127_c0 : nS_st4_b127_c1;
  assign nC_st5_b15_c0 = (nC_st4_b7_c0 == 0) ? nC_st4_b15_c0 : nC_st4_b15_c1;
  assign nC_st5_b31_c0 = (nC_st4_b23_c0 == 0) ? nC_st4_b31_c0 : nC_st4_b31_c1;
  assign nC_st5_b47_c0 = (nC_st4_b39_c0 == 0) ? nC_st4_b47_c0 : nC_st4_b47_c1;
  assign nC_st5_b63_c0 = (nC_st4_b55_c0 == 0) ? nC_st4_b63_c0 : nC_st4_b63_c1;
  assign nC_st5_b79_c0 = (nC_st4_b71_c0 == 0) ? nC_st4_b79_c0 : nC_st4_b79_c1;
  assign nC_st5_b95_c0 = (nC_st4_b87_c0 == 0) ? nC_st4_b95_c0 : nC_st4_b95_c1;
  assign nC_st5_b111_c0 = (nC_st4_b103_c0 == 0) ? nC_st4_b111_c0 : nC_st4_b111_c1;
  assign nC_st5_b127_c0 = (nC_st4_b119_c0 == 0) ? nC_st4_b127_c0 : nC_st4_b127_c1;
  assign nC_st5_b15_c1 = (nC_st4_b7_c1 == 0) ? nC_st4_b15_c0 : nC_st4_b15_c1;
  assign nC_st5_b31_c1 = (nC_st4_b23_c1 == 0) ? nC_st4_b31_c0 : nC_st4_b31_c1;
  assign nC_st5_b47_c1 = (nC_st4_b39_c1 == 0) ? nC_st4_b47_c0 : nC_st4_b47_c1;
  assign nC_st5_b63_c1 = (nC_st4_b55_c1 == 0) ? nC_st4_b63_c0 : nC_st4_b63_c1;
  assign nC_st5_b79_c1 = (nC_st4_b71_c1 == 0) ? nC_st4_b79_c0 : nC_st4_b79_c1;
  assign nC_st5_b95_c1 = (nC_st4_b87_c1 == 0) ? nC_st4_b95_c0 : nC_st4_b95_c1;
  assign nC_st5_b111_c1 = (nC_st4_b103_c1 == 0) ? nC_st4_b111_c0 : nC_st4_b111_c1;
  assign nC_st5_b127_c1 = (nC_st4_b119_c1 == 0) ? nC_st4_b127_c0 : nC_st4_b127_c1;

  assign nS_st6_b0_c0 = nS_st5_b0_c0;
  assign nS_st6_b1_c0 = nS_st5_b1_c0;
  assign nS_st6_b2_c0 = nS_st5_b2_c0;
  assign nS_st6_b3_c0 = nS_st5_b3_c0;
  assign nS_st6_b4_c0 = nS_st5_b4_c0;
  assign nS_st6_b5_c0 = nS_st5_b5_c0;
  assign nS_st6_b6_c0 = nS_st5_b6_c0;
  assign nS_st6_b7_c0 = nS_st5_b7_c0;
  assign nS_st6_b8_c0 = nS_st5_b8_c0;
  assign nS_st6_b9_c0 = nS_st5_b9_c0;
  assign nS_st6_b10_c0 = nS_st5_b10_c0;
  assign nS_st6_b11_c0 = nS_st5_b11_c0;
  assign nS_st6_b12_c0 = nS_st5_b12_c0;
  assign nS_st6_b13_c0 = nS_st5_b13_c0;
  assign nS_st6_b14_c0 = nS_st5_b14_c0;
  assign nS_st6_b15_c0 = nS_st5_b15_c0;
  assign nS_st6_b16_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b16_c0 : nS_st5_b16_c1;
  assign nS_st6_b17_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b17_c0 : nS_st5_b17_c1;
  assign nS_st6_b18_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b18_c0 : nS_st5_b18_c1;
  assign nS_st6_b19_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b19_c0 : nS_st5_b19_c1;
  assign nS_st6_b20_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b20_c0 : nS_st5_b20_c1;
  assign nS_st6_b21_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b21_c0 : nS_st5_b21_c1;
  assign nS_st6_b22_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b22_c0 : nS_st5_b22_c1;
  assign nS_st6_b23_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b23_c0 : nS_st5_b23_c1;
  assign nS_st6_b24_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b24_c0 : nS_st5_b24_c1;
  assign nS_st6_b25_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b25_c0 : nS_st5_b25_c1;
  assign nS_st6_b26_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b26_c0 : nS_st5_b26_c1;
  assign nS_st6_b27_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b27_c0 : nS_st5_b27_c1;
  assign nS_st6_b28_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b28_c0 : nS_st5_b28_c1;
  assign nS_st6_b29_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b29_c0 : nS_st5_b29_c1;
  assign nS_st6_b30_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b30_c0 : nS_st5_b30_c1;
  assign nS_st6_b31_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b31_c0 : nS_st5_b31_c1;
  assign nS_st6_b32_c0 = nS_st5_b32_c0;
  assign nS_st6_b33_c0 = nS_st5_b33_c0;
  assign nS_st6_b34_c0 = nS_st5_b34_c0;
  assign nS_st6_b35_c0 = nS_st5_b35_c0;
  assign nS_st6_b36_c0 = nS_st5_b36_c0;
  assign nS_st6_b37_c0 = nS_st5_b37_c0;
  assign nS_st6_b38_c0 = nS_st5_b38_c0;
  assign nS_st6_b39_c0 = nS_st5_b39_c0;
  assign nS_st6_b40_c0 = nS_st5_b40_c0;
  assign nS_st6_b41_c0 = nS_st5_b41_c0;
  assign nS_st6_b42_c0 = nS_st5_b42_c0;
  assign nS_st6_b43_c0 = nS_st5_b43_c0;
  assign nS_st6_b44_c0 = nS_st5_b44_c0;
  assign nS_st6_b45_c0 = nS_st5_b45_c0;
  assign nS_st6_b46_c0 = nS_st5_b46_c0;
  assign nS_st6_b47_c0 = nS_st5_b47_c0;
  assign nS_st6_b48_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b48_c0 : nS_st5_b48_c1;
  assign nS_st6_b49_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b49_c0 : nS_st5_b49_c1;
  assign nS_st6_b50_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b50_c0 : nS_st5_b50_c1;
  assign nS_st6_b51_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b51_c0 : nS_st5_b51_c1;
  assign nS_st6_b52_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b52_c0 : nS_st5_b52_c1;
  assign nS_st6_b53_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b53_c0 : nS_st5_b53_c1;
  assign nS_st6_b54_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b54_c0 : nS_st5_b54_c1;
  assign nS_st6_b55_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b55_c0 : nS_st5_b55_c1;
  assign nS_st6_b56_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b56_c0 : nS_st5_b56_c1;
  assign nS_st6_b57_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b57_c0 : nS_st5_b57_c1;
  assign nS_st6_b58_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b58_c0 : nS_st5_b58_c1;
  assign nS_st6_b59_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b59_c0 : nS_st5_b59_c1;
  assign nS_st6_b60_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b60_c0 : nS_st5_b60_c1;
  assign nS_st6_b61_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b61_c0 : nS_st5_b61_c1;
  assign nS_st6_b62_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b62_c0 : nS_st5_b62_c1;
  assign nS_st6_b63_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b63_c0 : nS_st5_b63_c1;
  assign nS_st6_b64_c0 = nS_st5_b64_c0;
  assign nS_st6_b65_c0 = nS_st5_b65_c0;
  assign nS_st6_b66_c0 = nS_st5_b66_c0;
  assign nS_st6_b67_c0 = nS_st5_b67_c0;
  assign nS_st6_b68_c0 = nS_st5_b68_c0;
  assign nS_st6_b69_c0 = nS_st5_b69_c0;
  assign nS_st6_b70_c0 = nS_st5_b70_c0;
  assign nS_st6_b71_c0 = nS_st5_b71_c0;
  assign nS_st6_b72_c0 = nS_st5_b72_c0;
  assign nS_st6_b73_c0 = nS_st5_b73_c0;
  assign nS_st6_b74_c0 = nS_st5_b74_c0;
  assign nS_st6_b75_c0 = nS_st5_b75_c0;
  assign nS_st6_b76_c0 = nS_st5_b76_c0;
  assign nS_st6_b77_c0 = nS_st5_b77_c0;
  assign nS_st6_b78_c0 = nS_st5_b78_c0;
  assign nS_st6_b79_c0 = nS_st5_b79_c0;
  assign nS_st6_b80_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b80_c0 : nS_st5_b80_c1;
  assign nS_st6_b81_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b81_c0 : nS_st5_b81_c1;
  assign nS_st6_b82_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b82_c0 : nS_st5_b82_c1;
  assign nS_st6_b83_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b83_c0 : nS_st5_b83_c1;
  assign nS_st6_b84_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b84_c0 : nS_st5_b84_c1;
  assign nS_st6_b85_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b85_c0 : nS_st5_b85_c1;
  assign nS_st6_b86_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b86_c0 : nS_st5_b86_c1;
  assign nS_st6_b87_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b87_c0 : nS_st5_b87_c1;
  assign nS_st6_b88_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b88_c0 : nS_st5_b88_c1;
  assign nS_st6_b89_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b89_c0 : nS_st5_b89_c1;
  assign nS_st6_b90_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b90_c0 : nS_st5_b90_c1;
  assign nS_st6_b91_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b91_c0 : nS_st5_b91_c1;
  assign nS_st6_b92_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b92_c0 : nS_st5_b92_c1;
  assign nS_st6_b93_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b93_c0 : nS_st5_b93_c1;
  assign nS_st6_b94_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b94_c0 : nS_st5_b94_c1;
  assign nS_st6_b95_c0 = (nC_st5_b79_c0 == 0) ? nS_st5_b95_c0 : nS_st5_b95_c1;
  assign nS_st6_b96_c0 = nS_st5_b96_c0;
  assign nS_st6_b97_c0 = nS_st5_b97_c0;
  assign nS_st6_b98_c0 = nS_st5_b98_c0;
  assign nS_st6_b99_c0 = nS_st5_b99_c0;
  assign nS_st6_b100_c0 = nS_st5_b100_c0;
  assign nS_st6_b101_c0 = nS_st5_b101_c0;
  assign nS_st6_b102_c0 = nS_st5_b102_c0;
  assign nS_st6_b103_c0 = nS_st5_b103_c0;
  assign nS_st6_b104_c0 = nS_st5_b104_c0;
  assign nS_st6_b105_c0 = nS_st5_b105_c0;
  assign nS_st6_b106_c0 = nS_st5_b106_c0;
  assign nS_st6_b107_c0 = nS_st5_b107_c0;
  assign nS_st6_b108_c0 = nS_st5_b108_c0;
  assign nS_st6_b109_c0 = nS_st5_b109_c0;
  assign nS_st6_b110_c0 = nS_st5_b110_c0;
  assign nS_st6_b111_c0 = nS_st5_b111_c0;
  assign nS_st6_b112_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b112_c0 : nS_st5_b112_c1;
  assign nS_st6_b113_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b113_c0 : nS_st5_b113_c1;
  assign nS_st6_b114_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b114_c0 : nS_st5_b114_c1;
  assign nS_st6_b115_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b115_c0 : nS_st5_b115_c1;
  assign nS_st6_b116_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b116_c0 : nS_st5_b116_c1;
  assign nS_st6_b117_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b117_c0 : nS_st5_b117_c1;
  assign nS_st6_b118_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b118_c0 : nS_st5_b118_c1;
  assign nS_st6_b119_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b119_c0 : nS_st5_b119_c1;
  assign nS_st6_b120_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b120_c0 : nS_st5_b120_c1;
  assign nS_st6_b121_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b121_c0 : nS_st5_b121_c1;
  assign nS_st6_b122_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b122_c0 : nS_st5_b122_c1;
  assign nS_st6_b123_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b123_c0 : nS_st5_b123_c1;
  assign nS_st6_b124_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b124_c0 : nS_st5_b124_c1;
  assign nS_st6_b125_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b125_c0 : nS_st5_b125_c1;
  assign nS_st6_b126_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b126_c0 : nS_st5_b126_c1;
  assign nS_st6_b127_c0 = (nC_st5_b111_c0 == 0) ? nS_st5_b127_c0 : nS_st5_b127_c1;
  assign nS_st6_b0_c1 = nS_st5_b0_c1;
  assign nS_st6_b1_c1 = nS_st5_b1_c1;
  assign nS_st6_b2_c1 = nS_st5_b2_c1;
  assign nS_st6_b3_c1 = nS_st5_b3_c1;
  assign nS_st6_b4_c1 = nS_st5_b4_c1;
  assign nS_st6_b5_c1 = nS_st5_b5_c1;
  assign nS_st6_b6_c1 = nS_st5_b6_c1;
  assign nS_st6_b7_c1 = nS_st5_b7_c1;
  assign nS_st6_b8_c1 = nS_st5_b8_c1;
  assign nS_st6_b9_c1 = nS_st5_b9_c1;
  assign nS_st6_b10_c1 = nS_st5_b10_c1;
  assign nS_st6_b11_c1 = nS_st5_b11_c1;
  assign nS_st6_b12_c1 = nS_st5_b12_c1;
  assign nS_st6_b13_c1 = nS_st5_b13_c1;
  assign nS_st6_b14_c1 = nS_st5_b14_c1;
  assign nS_st6_b15_c1 = nS_st5_b15_c1;
  assign nS_st6_b16_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b16_c0 : nS_st5_b16_c1;
  assign nS_st6_b17_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b17_c0 : nS_st5_b17_c1;
  assign nS_st6_b18_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b18_c0 : nS_st5_b18_c1;
  assign nS_st6_b19_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b19_c0 : nS_st5_b19_c1;
  assign nS_st6_b20_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b20_c0 : nS_st5_b20_c1;
  assign nS_st6_b21_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b21_c0 : nS_st5_b21_c1;
  assign nS_st6_b22_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b22_c0 : nS_st5_b22_c1;
  assign nS_st6_b23_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b23_c0 : nS_st5_b23_c1;
  assign nS_st6_b24_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b24_c0 : nS_st5_b24_c1;
  assign nS_st6_b25_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b25_c0 : nS_st5_b25_c1;
  assign nS_st6_b26_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b26_c0 : nS_st5_b26_c1;
  assign nS_st6_b27_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b27_c0 : nS_st5_b27_c1;
  assign nS_st6_b28_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b28_c0 : nS_st5_b28_c1;
  assign nS_st6_b29_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b29_c0 : nS_st5_b29_c1;
  assign nS_st6_b30_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b30_c0 : nS_st5_b30_c1;
  assign nS_st6_b31_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b31_c0 : nS_st5_b31_c1;
  assign nS_st6_b32_c1 = nS_st5_b32_c1;
  assign nS_st6_b33_c1 = nS_st5_b33_c1;
  assign nS_st6_b34_c1 = nS_st5_b34_c1;
  assign nS_st6_b35_c1 = nS_st5_b35_c1;
  assign nS_st6_b36_c1 = nS_st5_b36_c1;
  assign nS_st6_b37_c1 = nS_st5_b37_c1;
  assign nS_st6_b38_c1 = nS_st5_b38_c1;
  assign nS_st6_b39_c1 = nS_st5_b39_c1;
  assign nS_st6_b40_c1 = nS_st5_b40_c1;
  assign nS_st6_b41_c1 = nS_st5_b41_c1;
  assign nS_st6_b42_c1 = nS_st5_b42_c1;
  assign nS_st6_b43_c1 = nS_st5_b43_c1;
  assign nS_st6_b44_c1 = nS_st5_b44_c1;
  assign nS_st6_b45_c1 = nS_st5_b45_c1;
  assign nS_st6_b46_c1 = nS_st5_b46_c1;
  assign nS_st6_b47_c1 = nS_st5_b47_c1;
  assign nS_st6_b48_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b48_c0 : nS_st5_b48_c1;
  assign nS_st6_b49_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b49_c0 : nS_st5_b49_c1;
  assign nS_st6_b50_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b50_c0 : nS_st5_b50_c1;
  assign nS_st6_b51_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b51_c0 : nS_st5_b51_c1;
  assign nS_st6_b52_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b52_c0 : nS_st5_b52_c1;
  assign nS_st6_b53_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b53_c0 : nS_st5_b53_c1;
  assign nS_st6_b54_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b54_c0 : nS_st5_b54_c1;
  assign nS_st6_b55_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b55_c0 : nS_st5_b55_c1;
  assign nS_st6_b56_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b56_c0 : nS_st5_b56_c1;
  assign nS_st6_b57_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b57_c0 : nS_st5_b57_c1;
  assign nS_st6_b58_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b58_c0 : nS_st5_b58_c1;
  assign nS_st6_b59_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b59_c0 : nS_st5_b59_c1;
  assign nS_st6_b60_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b60_c0 : nS_st5_b60_c1;
  assign nS_st6_b61_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b61_c0 : nS_st5_b61_c1;
  assign nS_st6_b62_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b62_c0 : nS_st5_b62_c1;
  assign nS_st6_b63_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b63_c0 : nS_st5_b63_c1;
  assign nS_st6_b64_c1 = nS_st5_b64_c1;
  assign nS_st6_b65_c1 = nS_st5_b65_c1;
  assign nS_st6_b66_c1 = nS_st5_b66_c1;
  assign nS_st6_b67_c1 = nS_st5_b67_c1;
  assign nS_st6_b68_c1 = nS_st5_b68_c1;
  assign nS_st6_b69_c1 = nS_st5_b69_c1;
  assign nS_st6_b70_c1 = nS_st5_b70_c1;
  assign nS_st6_b71_c1 = nS_st5_b71_c1;
  assign nS_st6_b72_c1 = nS_st5_b72_c1;
  assign nS_st6_b73_c1 = nS_st5_b73_c1;
  assign nS_st6_b74_c1 = nS_st5_b74_c1;
  assign nS_st6_b75_c1 = nS_st5_b75_c1;
  assign nS_st6_b76_c1 = nS_st5_b76_c1;
  assign nS_st6_b77_c1 = nS_st5_b77_c1;
  assign nS_st6_b78_c1 = nS_st5_b78_c1;
  assign nS_st6_b79_c1 = nS_st5_b79_c1;
  assign nS_st6_b80_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b80_c0 : nS_st5_b80_c1;
  assign nS_st6_b81_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b81_c0 : nS_st5_b81_c1;
  assign nS_st6_b82_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b82_c0 : nS_st5_b82_c1;
  assign nS_st6_b83_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b83_c0 : nS_st5_b83_c1;
  assign nS_st6_b84_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b84_c0 : nS_st5_b84_c1;
  assign nS_st6_b85_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b85_c0 : nS_st5_b85_c1;
  assign nS_st6_b86_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b86_c0 : nS_st5_b86_c1;
  assign nS_st6_b87_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b87_c0 : nS_st5_b87_c1;
  assign nS_st6_b88_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b88_c0 : nS_st5_b88_c1;
  assign nS_st6_b89_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b89_c0 : nS_st5_b89_c1;
  assign nS_st6_b90_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b90_c0 : nS_st5_b90_c1;
  assign nS_st6_b91_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b91_c0 : nS_st5_b91_c1;
  assign nS_st6_b92_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b92_c0 : nS_st5_b92_c1;
  assign nS_st6_b93_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b93_c0 : nS_st5_b93_c1;
  assign nS_st6_b94_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b94_c0 : nS_st5_b94_c1;
  assign nS_st6_b95_c1 = (nC_st5_b79_c1 == 0) ? nS_st5_b95_c0 : nS_st5_b95_c1;
  assign nS_st6_b96_c1 = nS_st5_b96_c1;
  assign nS_st6_b97_c1 = nS_st5_b97_c1;
  assign nS_st6_b98_c1 = nS_st5_b98_c1;
  assign nS_st6_b99_c1 = nS_st5_b99_c1;
  assign nS_st6_b100_c1 = nS_st5_b100_c1;
  assign nS_st6_b101_c1 = nS_st5_b101_c1;
  assign nS_st6_b102_c1 = nS_st5_b102_c1;
  assign nS_st6_b103_c1 = nS_st5_b103_c1;
  assign nS_st6_b104_c1 = nS_st5_b104_c1;
  assign nS_st6_b105_c1 = nS_st5_b105_c1;
  assign nS_st6_b106_c1 = nS_st5_b106_c1;
  assign nS_st6_b107_c1 = nS_st5_b107_c1;
  assign nS_st6_b108_c1 = nS_st5_b108_c1;
  assign nS_st6_b109_c1 = nS_st5_b109_c1;
  assign nS_st6_b110_c1 = nS_st5_b110_c1;
  assign nS_st6_b111_c1 = nS_st5_b111_c1;
  assign nS_st6_b112_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b112_c0 : nS_st5_b112_c1;
  assign nS_st6_b113_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b113_c0 : nS_st5_b113_c1;
  assign nS_st6_b114_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b114_c0 : nS_st5_b114_c1;
  assign nS_st6_b115_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b115_c0 : nS_st5_b115_c1;
  assign nS_st6_b116_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b116_c0 : nS_st5_b116_c1;
  assign nS_st6_b117_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b117_c0 : nS_st5_b117_c1;
  assign nS_st6_b118_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b118_c0 : nS_st5_b118_c1;
  assign nS_st6_b119_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b119_c0 : nS_st5_b119_c1;
  assign nS_st6_b120_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b120_c0 : nS_st5_b120_c1;
  assign nS_st6_b121_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b121_c0 : nS_st5_b121_c1;
  assign nS_st6_b122_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b122_c0 : nS_st5_b122_c1;
  assign nS_st6_b123_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b123_c0 : nS_st5_b123_c1;
  assign nS_st6_b124_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b124_c0 : nS_st5_b124_c1;
  assign nS_st6_b125_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b125_c0 : nS_st5_b125_c1;
  assign nS_st6_b126_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b126_c0 : nS_st5_b126_c1;
  assign nS_st6_b127_c1 = (nC_st5_b111_c1 == 0) ? nS_st5_b127_c0 : nS_st5_b127_c1;
  assign nC_st6_b31_c0 = (nC_st5_b15_c0 == 0) ? nC_st5_b31_c0 : nC_st5_b31_c1;
  assign nC_st6_b63_c0 = (nC_st5_b47_c0 == 0) ? nC_st5_b63_c0 : nC_st5_b63_c1;
  assign nC_st6_b95_c0 = (nC_st5_b79_c0 == 0) ? nC_st5_b95_c0 : nC_st5_b95_c1;
  assign nC_st6_b127_c0 = (nC_st5_b111_c0 == 0) ? nC_st5_b127_c0 : nC_st5_b127_c1;
  assign nC_st6_b31_c1 = (nC_st5_b15_c1 == 0) ? nC_st5_b31_c0 : nC_st5_b31_c1;
  assign nC_st6_b63_c1 = (nC_st5_b47_c1 == 0) ? nC_st5_b63_c0 : nC_st5_b63_c1;
  assign nC_st6_b95_c1 = (nC_st5_b79_c1 == 0) ? nC_st5_b95_c0 : nC_st5_b95_c1;
  assign nC_st6_b127_c1 = (nC_st5_b111_c1 == 0) ? nC_st5_b127_c0 : nC_st5_b127_c1;

  assign nS_st7_b0_c0 = nS_st6_b0_c0;
  assign nS_st7_b1_c0 = nS_st6_b1_c0;
  assign nS_st7_b2_c0 = nS_st6_b2_c0;
  assign nS_st7_b3_c0 = nS_st6_b3_c0;
  assign nS_st7_b4_c0 = nS_st6_b4_c0;
  assign nS_st7_b5_c0 = nS_st6_b5_c0;
  assign nS_st7_b6_c0 = nS_st6_b6_c0;
  assign nS_st7_b7_c0 = nS_st6_b7_c0;
  assign nS_st7_b8_c0 = nS_st6_b8_c0;
  assign nS_st7_b9_c0 = nS_st6_b9_c0;
  assign nS_st7_b10_c0 = nS_st6_b10_c0;
  assign nS_st7_b11_c0 = nS_st6_b11_c0;
  assign nS_st7_b12_c0 = nS_st6_b12_c0;
  assign nS_st7_b13_c0 = nS_st6_b13_c0;
  assign nS_st7_b14_c0 = nS_st6_b14_c0;
  assign nS_st7_b15_c0 = nS_st6_b15_c0;
  assign nS_st7_b16_c0 = nS_st6_b16_c0;
  assign nS_st7_b17_c0 = nS_st6_b17_c0;
  assign nS_st7_b18_c0 = nS_st6_b18_c0;
  assign nS_st7_b19_c0 = nS_st6_b19_c0;
  assign nS_st7_b20_c0 = nS_st6_b20_c0;
  assign nS_st7_b21_c0 = nS_st6_b21_c0;
  assign nS_st7_b22_c0 = nS_st6_b22_c0;
  assign nS_st7_b23_c0 = nS_st6_b23_c0;
  assign nS_st7_b24_c0 = nS_st6_b24_c0;
  assign nS_st7_b25_c0 = nS_st6_b25_c0;
  assign nS_st7_b26_c0 = nS_st6_b26_c0;
  assign nS_st7_b27_c0 = nS_st6_b27_c0;
  assign nS_st7_b28_c0 = nS_st6_b28_c0;
  assign nS_st7_b29_c0 = nS_st6_b29_c0;
  assign nS_st7_b30_c0 = nS_st6_b30_c0;
  assign nS_st7_b31_c0 = nS_st6_b31_c0;
  assign nS_st7_b32_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b32_c0 : nS_st6_b32_c1;
  assign nS_st7_b33_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b33_c0 : nS_st6_b33_c1;
  assign nS_st7_b34_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b34_c0 : nS_st6_b34_c1;
  assign nS_st7_b35_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b35_c0 : nS_st6_b35_c1;
  assign nS_st7_b36_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b36_c0 : nS_st6_b36_c1;
  assign nS_st7_b37_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b37_c0 : nS_st6_b37_c1;
  assign nS_st7_b38_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b38_c0 : nS_st6_b38_c1;
  assign nS_st7_b39_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b39_c0 : nS_st6_b39_c1;
  assign nS_st7_b40_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b40_c0 : nS_st6_b40_c1;
  assign nS_st7_b41_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b41_c0 : nS_st6_b41_c1;
  assign nS_st7_b42_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b42_c0 : nS_st6_b42_c1;
  assign nS_st7_b43_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b43_c0 : nS_st6_b43_c1;
  assign nS_st7_b44_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b44_c0 : nS_st6_b44_c1;
  assign nS_st7_b45_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b45_c0 : nS_st6_b45_c1;
  assign nS_st7_b46_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b46_c0 : nS_st6_b46_c1;
  assign nS_st7_b47_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b47_c0 : nS_st6_b47_c1;
  assign nS_st7_b48_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b48_c0 : nS_st6_b48_c1;
  assign nS_st7_b49_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b49_c0 : nS_st6_b49_c1;
  assign nS_st7_b50_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b50_c0 : nS_st6_b50_c1;
  assign nS_st7_b51_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b51_c0 : nS_st6_b51_c1;
  assign nS_st7_b52_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b52_c0 : nS_st6_b52_c1;
  assign nS_st7_b53_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b53_c0 : nS_st6_b53_c1;
  assign nS_st7_b54_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b54_c0 : nS_st6_b54_c1;
  assign nS_st7_b55_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b55_c0 : nS_st6_b55_c1;
  assign nS_st7_b56_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b56_c0 : nS_st6_b56_c1;
  assign nS_st7_b57_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b57_c0 : nS_st6_b57_c1;
  assign nS_st7_b58_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b58_c0 : nS_st6_b58_c1;
  assign nS_st7_b59_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b59_c0 : nS_st6_b59_c1;
  assign nS_st7_b60_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b60_c0 : nS_st6_b60_c1;
  assign nS_st7_b61_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b61_c0 : nS_st6_b61_c1;
  assign nS_st7_b62_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b62_c0 : nS_st6_b62_c1;
  assign nS_st7_b63_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b63_c0 : nS_st6_b63_c1;
  assign nS_st7_b64_c0 = nS_st6_b64_c0;
  assign nS_st7_b65_c0 = nS_st6_b65_c0;
  assign nS_st7_b66_c0 = nS_st6_b66_c0;
  assign nS_st7_b67_c0 = nS_st6_b67_c0;
  assign nS_st7_b68_c0 = nS_st6_b68_c0;
  assign nS_st7_b69_c0 = nS_st6_b69_c0;
  assign nS_st7_b70_c0 = nS_st6_b70_c0;
  assign nS_st7_b71_c0 = nS_st6_b71_c0;
  assign nS_st7_b72_c0 = nS_st6_b72_c0;
  assign nS_st7_b73_c0 = nS_st6_b73_c0;
  assign nS_st7_b74_c0 = nS_st6_b74_c0;
  assign nS_st7_b75_c0 = nS_st6_b75_c0;
  assign nS_st7_b76_c0 = nS_st6_b76_c0;
  assign nS_st7_b77_c0 = nS_st6_b77_c0;
  assign nS_st7_b78_c0 = nS_st6_b78_c0;
  assign nS_st7_b79_c0 = nS_st6_b79_c0;
  assign nS_st7_b80_c0 = nS_st6_b80_c0;
  assign nS_st7_b81_c0 = nS_st6_b81_c0;
  assign nS_st7_b82_c0 = nS_st6_b82_c0;
  assign nS_st7_b83_c0 = nS_st6_b83_c0;
  assign nS_st7_b84_c0 = nS_st6_b84_c0;
  assign nS_st7_b85_c0 = nS_st6_b85_c0;
  assign nS_st7_b86_c0 = nS_st6_b86_c0;
  assign nS_st7_b87_c0 = nS_st6_b87_c0;
  assign nS_st7_b88_c0 = nS_st6_b88_c0;
  assign nS_st7_b89_c0 = nS_st6_b89_c0;
  assign nS_st7_b90_c0 = nS_st6_b90_c0;
  assign nS_st7_b91_c0 = nS_st6_b91_c0;
  assign nS_st7_b92_c0 = nS_st6_b92_c0;
  assign nS_st7_b93_c0 = nS_st6_b93_c0;
  assign nS_st7_b94_c0 = nS_st6_b94_c0;
  assign nS_st7_b95_c0 = nS_st6_b95_c0;
  assign nS_st7_b96_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b96_c0 : nS_st6_b96_c1;
  assign nS_st7_b97_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b97_c0 : nS_st6_b97_c1;
  assign nS_st7_b98_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b98_c0 : nS_st6_b98_c1;
  assign nS_st7_b99_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b99_c0 : nS_st6_b99_c1;
  assign nS_st7_b100_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b100_c0 : nS_st6_b100_c1;
  assign nS_st7_b101_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b101_c0 : nS_st6_b101_c1;
  assign nS_st7_b102_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b102_c0 : nS_st6_b102_c1;
  assign nS_st7_b103_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b103_c0 : nS_st6_b103_c1;
  assign nS_st7_b104_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b104_c0 : nS_st6_b104_c1;
  assign nS_st7_b105_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b105_c0 : nS_st6_b105_c1;
  assign nS_st7_b106_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b106_c0 : nS_st6_b106_c1;
  assign nS_st7_b107_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b107_c0 : nS_st6_b107_c1;
  assign nS_st7_b108_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b108_c0 : nS_st6_b108_c1;
  assign nS_st7_b109_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b109_c0 : nS_st6_b109_c1;
  assign nS_st7_b110_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b110_c0 : nS_st6_b110_c1;
  assign nS_st7_b111_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b111_c0 : nS_st6_b111_c1;
  assign nS_st7_b112_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b112_c0 : nS_st6_b112_c1;
  assign nS_st7_b113_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b113_c0 : nS_st6_b113_c1;
  assign nS_st7_b114_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b114_c0 : nS_st6_b114_c1;
  assign nS_st7_b115_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b115_c0 : nS_st6_b115_c1;
  assign nS_st7_b116_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b116_c0 : nS_st6_b116_c1;
  assign nS_st7_b117_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b117_c0 : nS_st6_b117_c1;
  assign nS_st7_b118_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b118_c0 : nS_st6_b118_c1;
  assign nS_st7_b119_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b119_c0 : nS_st6_b119_c1;
  assign nS_st7_b120_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b120_c0 : nS_st6_b120_c1;
  assign nS_st7_b121_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b121_c0 : nS_st6_b121_c1;
  assign nS_st7_b122_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b122_c0 : nS_st6_b122_c1;
  assign nS_st7_b123_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b123_c0 : nS_st6_b123_c1;
  assign nS_st7_b124_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b124_c0 : nS_st6_b124_c1;
  assign nS_st7_b125_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b125_c0 : nS_st6_b125_c1;
  assign nS_st7_b126_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b126_c0 : nS_st6_b126_c1;
  assign nS_st7_b127_c0 = (nC_st6_b95_c0 == 0) ? nS_st6_b127_c0 : nS_st6_b127_c1;
  assign nS_st7_b0_c1 = nS_st6_b0_c1;
  assign nS_st7_b1_c1 = nS_st6_b1_c1;
  assign nS_st7_b2_c1 = nS_st6_b2_c1;
  assign nS_st7_b3_c1 = nS_st6_b3_c1;
  assign nS_st7_b4_c1 = nS_st6_b4_c1;
  assign nS_st7_b5_c1 = nS_st6_b5_c1;
  assign nS_st7_b6_c1 = nS_st6_b6_c1;
  assign nS_st7_b7_c1 = nS_st6_b7_c1;
  assign nS_st7_b8_c1 = nS_st6_b8_c1;
  assign nS_st7_b9_c1 = nS_st6_b9_c1;
  assign nS_st7_b10_c1 = nS_st6_b10_c1;
  assign nS_st7_b11_c1 = nS_st6_b11_c1;
  assign nS_st7_b12_c1 = nS_st6_b12_c1;
  assign nS_st7_b13_c1 = nS_st6_b13_c1;
  assign nS_st7_b14_c1 = nS_st6_b14_c1;
  assign nS_st7_b15_c1 = nS_st6_b15_c1;
  assign nS_st7_b16_c1 = nS_st6_b16_c1;
  assign nS_st7_b17_c1 = nS_st6_b17_c1;
  assign nS_st7_b18_c1 = nS_st6_b18_c1;
  assign nS_st7_b19_c1 = nS_st6_b19_c1;
  assign nS_st7_b20_c1 = nS_st6_b20_c1;
  assign nS_st7_b21_c1 = nS_st6_b21_c1;
  assign nS_st7_b22_c1 = nS_st6_b22_c1;
  assign nS_st7_b23_c1 = nS_st6_b23_c1;
  assign nS_st7_b24_c1 = nS_st6_b24_c1;
  assign nS_st7_b25_c1 = nS_st6_b25_c1;
  assign nS_st7_b26_c1 = nS_st6_b26_c1;
  assign nS_st7_b27_c1 = nS_st6_b27_c1;
  assign nS_st7_b28_c1 = nS_st6_b28_c1;
  assign nS_st7_b29_c1 = nS_st6_b29_c1;
  assign nS_st7_b30_c1 = nS_st6_b30_c1;
  assign nS_st7_b31_c1 = nS_st6_b31_c1;
  assign nS_st7_b32_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b32_c0 : nS_st6_b32_c1;
  assign nS_st7_b33_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b33_c0 : nS_st6_b33_c1;
  assign nS_st7_b34_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b34_c0 : nS_st6_b34_c1;
  assign nS_st7_b35_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b35_c0 : nS_st6_b35_c1;
  assign nS_st7_b36_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b36_c0 : nS_st6_b36_c1;
  assign nS_st7_b37_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b37_c0 : nS_st6_b37_c1;
  assign nS_st7_b38_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b38_c0 : nS_st6_b38_c1;
  assign nS_st7_b39_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b39_c0 : nS_st6_b39_c1;
  assign nS_st7_b40_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b40_c0 : nS_st6_b40_c1;
  assign nS_st7_b41_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b41_c0 : nS_st6_b41_c1;
  assign nS_st7_b42_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b42_c0 : nS_st6_b42_c1;
  assign nS_st7_b43_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b43_c0 : nS_st6_b43_c1;
  assign nS_st7_b44_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b44_c0 : nS_st6_b44_c1;
  assign nS_st7_b45_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b45_c0 : nS_st6_b45_c1;
  assign nS_st7_b46_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b46_c0 : nS_st6_b46_c1;
  assign nS_st7_b47_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b47_c0 : nS_st6_b47_c1;
  assign nS_st7_b48_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b48_c0 : nS_st6_b48_c1;
  assign nS_st7_b49_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b49_c0 : nS_st6_b49_c1;
  assign nS_st7_b50_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b50_c0 : nS_st6_b50_c1;
  assign nS_st7_b51_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b51_c0 : nS_st6_b51_c1;
  assign nS_st7_b52_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b52_c0 : nS_st6_b52_c1;
  assign nS_st7_b53_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b53_c0 : nS_st6_b53_c1;
  assign nS_st7_b54_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b54_c0 : nS_st6_b54_c1;
  assign nS_st7_b55_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b55_c0 : nS_st6_b55_c1;
  assign nS_st7_b56_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b56_c0 : nS_st6_b56_c1;
  assign nS_st7_b57_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b57_c0 : nS_st6_b57_c1;
  assign nS_st7_b58_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b58_c0 : nS_st6_b58_c1;
  assign nS_st7_b59_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b59_c0 : nS_st6_b59_c1;
  assign nS_st7_b60_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b60_c0 : nS_st6_b60_c1;
  assign nS_st7_b61_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b61_c0 : nS_st6_b61_c1;
  assign nS_st7_b62_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b62_c0 : nS_st6_b62_c1;
  assign nS_st7_b63_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b63_c0 : nS_st6_b63_c1;
  assign nS_st7_b64_c1 = nS_st6_b64_c1;
  assign nS_st7_b65_c1 = nS_st6_b65_c1;
  assign nS_st7_b66_c1 = nS_st6_b66_c1;
  assign nS_st7_b67_c1 = nS_st6_b67_c1;
  assign nS_st7_b68_c1 = nS_st6_b68_c1;
  assign nS_st7_b69_c1 = nS_st6_b69_c1;
  assign nS_st7_b70_c1 = nS_st6_b70_c1;
  assign nS_st7_b71_c1 = nS_st6_b71_c1;
  assign nS_st7_b72_c1 = nS_st6_b72_c1;
  assign nS_st7_b73_c1 = nS_st6_b73_c1;
  assign nS_st7_b74_c1 = nS_st6_b74_c1;
  assign nS_st7_b75_c1 = nS_st6_b75_c1;
  assign nS_st7_b76_c1 = nS_st6_b76_c1;
  assign nS_st7_b77_c1 = nS_st6_b77_c1;
  assign nS_st7_b78_c1 = nS_st6_b78_c1;
  assign nS_st7_b79_c1 = nS_st6_b79_c1;
  assign nS_st7_b80_c1 = nS_st6_b80_c1;
  assign nS_st7_b81_c1 = nS_st6_b81_c1;
  assign nS_st7_b82_c1 = nS_st6_b82_c1;
  assign nS_st7_b83_c1 = nS_st6_b83_c1;
  assign nS_st7_b84_c1 = nS_st6_b84_c1;
  assign nS_st7_b85_c1 = nS_st6_b85_c1;
  assign nS_st7_b86_c1 = nS_st6_b86_c1;
  assign nS_st7_b87_c1 = nS_st6_b87_c1;
  assign nS_st7_b88_c1 = nS_st6_b88_c1;
  assign nS_st7_b89_c1 = nS_st6_b89_c1;
  assign nS_st7_b90_c1 = nS_st6_b90_c1;
  assign nS_st7_b91_c1 = nS_st6_b91_c1;
  assign nS_st7_b92_c1 = nS_st6_b92_c1;
  assign nS_st7_b93_c1 = nS_st6_b93_c1;
  assign nS_st7_b94_c1 = nS_st6_b94_c1;
  assign nS_st7_b95_c1 = nS_st6_b95_c1;
  assign nS_st7_b96_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b96_c0 : nS_st6_b96_c1;
  assign nS_st7_b97_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b97_c0 : nS_st6_b97_c1;
  assign nS_st7_b98_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b98_c0 : nS_st6_b98_c1;
  assign nS_st7_b99_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b99_c0 : nS_st6_b99_c1;
  assign nS_st7_b100_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b100_c0 : nS_st6_b100_c1;
  assign nS_st7_b101_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b101_c0 : nS_st6_b101_c1;
  assign nS_st7_b102_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b102_c0 : nS_st6_b102_c1;
  assign nS_st7_b103_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b103_c0 : nS_st6_b103_c1;
  assign nS_st7_b104_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b104_c0 : nS_st6_b104_c1;
  assign nS_st7_b105_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b105_c0 : nS_st6_b105_c1;
  assign nS_st7_b106_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b106_c0 : nS_st6_b106_c1;
  assign nS_st7_b107_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b107_c0 : nS_st6_b107_c1;
  assign nS_st7_b108_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b108_c0 : nS_st6_b108_c1;
  assign nS_st7_b109_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b109_c0 : nS_st6_b109_c1;
  assign nS_st7_b110_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b110_c0 : nS_st6_b110_c1;
  assign nS_st7_b111_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b111_c0 : nS_st6_b111_c1;
  assign nS_st7_b112_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b112_c0 : nS_st6_b112_c1;
  assign nS_st7_b113_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b113_c0 : nS_st6_b113_c1;
  assign nS_st7_b114_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b114_c0 : nS_st6_b114_c1;
  assign nS_st7_b115_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b115_c0 : nS_st6_b115_c1;
  assign nS_st7_b116_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b116_c0 : nS_st6_b116_c1;
  assign nS_st7_b117_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b117_c0 : nS_st6_b117_c1;
  assign nS_st7_b118_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b118_c0 : nS_st6_b118_c1;
  assign nS_st7_b119_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b119_c0 : nS_st6_b119_c1;
  assign nS_st7_b120_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b120_c0 : nS_st6_b120_c1;
  assign nS_st7_b121_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b121_c0 : nS_st6_b121_c1;
  assign nS_st7_b122_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b122_c0 : nS_st6_b122_c1;
  assign nS_st7_b123_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b123_c0 : nS_st6_b123_c1;
  assign nS_st7_b124_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b124_c0 : nS_st6_b124_c1;
  assign nS_st7_b125_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b125_c0 : nS_st6_b125_c1;
  assign nS_st7_b126_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b126_c0 : nS_st6_b126_c1;
  assign nS_st7_b127_c1 = (nC_st6_b95_c1 == 0) ? nS_st6_b127_c0 : nS_st6_b127_c1;
  assign nC_st7_b63_c0 = (nC_st6_b31_c0 == 0) ? nC_st6_b63_c0 : nC_st6_b63_c1;
  assign nC_st7_b127_c0 = (nC_st6_b95_c0 == 0) ? nC_st6_b127_c0 : nC_st6_b127_c1;
  assign nC_st7_b63_c1 = (nC_st6_b31_c1 == 0) ? nC_st6_b63_c0 : nC_st6_b63_c1;
  assign nC_st7_b127_c1 = (nC_st6_b95_c1 == 0) ? nC_st6_b127_c0 : nC_st6_b127_c1;

  assign nS_st8_b0_c0 = nS_st7_b0_c0;
  assign nS_st8_b1_c0 = nS_st7_b1_c0;
  assign nS_st8_b2_c0 = nS_st7_b2_c0;
  assign nS_st8_b3_c0 = nS_st7_b3_c0;
  assign nS_st8_b4_c0 = nS_st7_b4_c0;
  assign nS_st8_b5_c0 = nS_st7_b5_c0;
  assign nS_st8_b6_c0 = nS_st7_b6_c0;
  assign nS_st8_b7_c0 = nS_st7_b7_c0;
  assign nS_st8_b8_c0 = nS_st7_b8_c0;
  assign nS_st8_b9_c0 = nS_st7_b9_c0;
  assign nS_st8_b10_c0 = nS_st7_b10_c0;
  assign nS_st8_b11_c0 = nS_st7_b11_c0;
  assign nS_st8_b12_c0 = nS_st7_b12_c0;
  assign nS_st8_b13_c0 = nS_st7_b13_c0;
  assign nS_st8_b14_c0 = nS_st7_b14_c0;
  assign nS_st8_b15_c0 = nS_st7_b15_c0;
  assign nS_st8_b16_c0 = nS_st7_b16_c0;
  assign nS_st8_b17_c0 = nS_st7_b17_c0;
  assign nS_st8_b18_c0 = nS_st7_b18_c0;
  assign nS_st8_b19_c0 = nS_st7_b19_c0;
  assign nS_st8_b20_c0 = nS_st7_b20_c0;
  assign nS_st8_b21_c0 = nS_st7_b21_c0;
  assign nS_st8_b22_c0 = nS_st7_b22_c0;
  assign nS_st8_b23_c0 = nS_st7_b23_c0;
  assign nS_st8_b24_c0 = nS_st7_b24_c0;
  assign nS_st8_b25_c0 = nS_st7_b25_c0;
  assign nS_st8_b26_c0 = nS_st7_b26_c0;
  assign nS_st8_b27_c0 = nS_st7_b27_c0;
  assign nS_st8_b28_c0 = nS_st7_b28_c0;
  assign nS_st8_b29_c0 = nS_st7_b29_c0;
  assign nS_st8_b30_c0 = nS_st7_b30_c0;
  assign nS_st8_b31_c0 = nS_st7_b31_c0;
  assign nS_st8_b32_c0 = nS_st7_b32_c0;
  assign nS_st8_b33_c0 = nS_st7_b33_c0;
  assign nS_st8_b34_c0 = nS_st7_b34_c0;
  assign nS_st8_b35_c0 = nS_st7_b35_c0;
  assign nS_st8_b36_c0 = nS_st7_b36_c0;
  assign nS_st8_b37_c0 = nS_st7_b37_c0;
  assign nS_st8_b38_c0 = nS_st7_b38_c0;
  assign nS_st8_b39_c0 = nS_st7_b39_c0;
  assign nS_st8_b40_c0 = nS_st7_b40_c0;
  assign nS_st8_b41_c0 = nS_st7_b41_c0;
  assign nS_st8_b42_c0 = nS_st7_b42_c0;
  assign nS_st8_b43_c0 = nS_st7_b43_c0;
  assign nS_st8_b44_c0 = nS_st7_b44_c0;
  assign nS_st8_b45_c0 = nS_st7_b45_c0;
  assign nS_st8_b46_c0 = nS_st7_b46_c0;
  assign nS_st8_b47_c0 = nS_st7_b47_c0;
  assign nS_st8_b48_c0 = nS_st7_b48_c0;
  assign nS_st8_b49_c0 = nS_st7_b49_c0;
  assign nS_st8_b50_c0 = nS_st7_b50_c0;
  assign nS_st8_b51_c0 = nS_st7_b51_c0;
  assign nS_st8_b52_c0 = nS_st7_b52_c0;
  assign nS_st8_b53_c0 = nS_st7_b53_c0;
  assign nS_st8_b54_c0 = nS_st7_b54_c0;
  assign nS_st8_b55_c0 = nS_st7_b55_c0;
  assign nS_st8_b56_c0 = nS_st7_b56_c0;
  assign nS_st8_b57_c0 = nS_st7_b57_c0;
  assign nS_st8_b58_c0 = nS_st7_b58_c0;
  assign nS_st8_b59_c0 = nS_st7_b59_c0;
  assign nS_st8_b60_c0 = nS_st7_b60_c0;
  assign nS_st8_b61_c0 = nS_st7_b61_c0;
  assign nS_st8_b62_c0 = nS_st7_b62_c0;
  assign nS_st8_b63_c0 = nS_st7_b63_c0;
  assign nS_st8_b64_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b64_c0 : nS_st7_b64_c1;
  assign nS_st8_b65_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b65_c0 : nS_st7_b65_c1;
  assign nS_st8_b66_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b66_c0 : nS_st7_b66_c1;
  assign nS_st8_b67_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b67_c0 : nS_st7_b67_c1;
  assign nS_st8_b68_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b68_c0 : nS_st7_b68_c1;
  assign nS_st8_b69_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b69_c0 : nS_st7_b69_c1;
  assign nS_st8_b70_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b70_c0 : nS_st7_b70_c1;
  assign nS_st8_b71_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b71_c0 : nS_st7_b71_c1;
  assign nS_st8_b72_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b72_c0 : nS_st7_b72_c1;
  assign nS_st8_b73_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b73_c0 : nS_st7_b73_c1;
  assign nS_st8_b74_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b74_c0 : nS_st7_b74_c1;
  assign nS_st8_b75_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b75_c0 : nS_st7_b75_c1;
  assign nS_st8_b76_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b76_c0 : nS_st7_b76_c1;
  assign nS_st8_b77_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b77_c0 : nS_st7_b77_c1;
  assign nS_st8_b78_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b78_c0 : nS_st7_b78_c1;
  assign nS_st8_b79_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b79_c0 : nS_st7_b79_c1;
  assign nS_st8_b80_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b80_c0 : nS_st7_b80_c1;
  assign nS_st8_b81_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b81_c0 : nS_st7_b81_c1;
  assign nS_st8_b82_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b82_c0 : nS_st7_b82_c1;
  assign nS_st8_b83_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b83_c0 : nS_st7_b83_c1;
  assign nS_st8_b84_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b84_c0 : nS_st7_b84_c1;
  assign nS_st8_b85_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b85_c0 : nS_st7_b85_c1;
  assign nS_st8_b86_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b86_c0 : nS_st7_b86_c1;
  assign nS_st8_b87_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b87_c0 : nS_st7_b87_c1;
  assign nS_st8_b88_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b88_c0 : nS_st7_b88_c1;
  assign nS_st8_b89_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b89_c0 : nS_st7_b89_c1;
  assign nS_st8_b90_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b90_c0 : nS_st7_b90_c1;
  assign nS_st8_b91_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b91_c0 : nS_st7_b91_c1;
  assign nS_st8_b92_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b92_c0 : nS_st7_b92_c1;
  assign nS_st8_b93_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b93_c0 : nS_st7_b93_c1;
  assign nS_st8_b94_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b94_c0 : nS_st7_b94_c1;
  assign nS_st8_b95_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b95_c0 : nS_st7_b95_c1;
  assign nS_st8_b96_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b96_c0 : nS_st7_b96_c1;
  assign nS_st8_b97_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b97_c0 : nS_st7_b97_c1;
  assign nS_st8_b98_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b98_c0 : nS_st7_b98_c1;
  assign nS_st8_b99_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b99_c0 : nS_st7_b99_c1;
  assign nS_st8_b100_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b100_c0 : nS_st7_b100_c1;
  assign nS_st8_b101_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b101_c0 : nS_st7_b101_c1;
  assign nS_st8_b102_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b102_c0 : nS_st7_b102_c1;
  assign nS_st8_b103_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b103_c0 : nS_st7_b103_c1;
  assign nS_st8_b104_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b104_c0 : nS_st7_b104_c1;
  assign nS_st8_b105_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b105_c0 : nS_st7_b105_c1;
  assign nS_st8_b106_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b106_c0 : nS_st7_b106_c1;
  assign nS_st8_b107_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b107_c0 : nS_st7_b107_c1;
  assign nS_st8_b108_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b108_c0 : nS_st7_b108_c1;
  assign nS_st8_b109_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b109_c0 : nS_st7_b109_c1;
  assign nS_st8_b110_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b110_c0 : nS_st7_b110_c1;
  assign nS_st8_b111_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b111_c0 : nS_st7_b111_c1;
  assign nS_st8_b112_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b112_c0 : nS_st7_b112_c1;
  assign nS_st8_b113_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b113_c0 : nS_st7_b113_c1;
  assign nS_st8_b114_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b114_c0 : nS_st7_b114_c1;
  assign nS_st8_b115_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b115_c0 : nS_st7_b115_c1;
  assign nS_st8_b116_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b116_c0 : nS_st7_b116_c1;
  assign nS_st8_b117_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b117_c0 : nS_st7_b117_c1;
  assign nS_st8_b118_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b118_c0 : nS_st7_b118_c1;
  assign nS_st8_b119_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b119_c0 : nS_st7_b119_c1;
  assign nS_st8_b120_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b120_c0 : nS_st7_b120_c1;
  assign nS_st8_b121_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b121_c0 : nS_st7_b121_c1;
  assign nS_st8_b122_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b122_c0 : nS_st7_b122_c1;
  assign nS_st8_b123_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b123_c0 : nS_st7_b123_c1;
  assign nS_st8_b124_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b124_c0 : nS_st7_b124_c1;
  assign nS_st8_b125_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b125_c0 : nS_st7_b125_c1;
  assign nS_st8_b126_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b126_c0 : nS_st7_b126_c1;
  assign nS_st8_b127_c0 = (nC_st7_b63_c0 == 0) ? nS_st7_b127_c0 : nS_st7_b127_c1;
  assign nS_st8_b0_c1 = nS_st7_b0_c1;
  assign nS_st8_b1_c1 = nS_st7_b1_c1;
  assign nS_st8_b2_c1 = nS_st7_b2_c1;
  assign nS_st8_b3_c1 = nS_st7_b3_c1;
  assign nS_st8_b4_c1 = nS_st7_b4_c1;
  assign nS_st8_b5_c1 = nS_st7_b5_c1;
  assign nS_st8_b6_c1 = nS_st7_b6_c1;
  assign nS_st8_b7_c1 = nS_st7_b7_c1;
  assign nS_st8_b8_c1 = nS_st7_b8_c1;
  assign nS_st8_b9_c1 = nS_st7_b9_c1;
  assign nS_st8_b10_c1 = nS_st7_b10_c1;
  assign nS_st8_b11_c1 = nS_st7_b11_c1;
  assign nS_st8_b12_c1 = nS_st7_b12_c1;
  assign nS_st8_b13_c1 = nS_st7_b13_c1;
  assign nS_st8_b14_c1 = nS_st7_b14_c1;
  assign nS_st8_b15_c1 = nS_st7_b15_c1;
  assign nS_st8_b16_c1 = nS_st7_b16_c1;
  assign nS_st8_b17_c1 = nS_st7_b17_c1;
  assign nS_st8_b18_c1 = nS_st7_b18_c1;
  assign nS_st8_b19_c1 = nS_st7_b19_c1;
  assign nS_st8_b20_c1 = nS_st7_b20_c1;
  assign nS_st8_b21_c1 = nS_st7_b21_c1;
  assign nS_st8_b22_c1 = nS_st7_b22_c1;
  assign nS_st8_b23_c1 = nS_st7_b23_c1;
  assign nS_st8_b24_c1 = nS_st7_b24_c1;
  assign nS_st8_b25_c1 = nS_st7_b25_c1;
  assign nS_st8_b26_c1 = nS_st7_b26_c1;
  assign nS_st8_b27_c1 = nS_st7_b27_c1;
  assign nS_st8_b28_c1 = nS_st7_b28_c1;
  assign nS_st8_b29_c1 = nS_st7_b29_c1;
  assign nS_st8_b30_c1 = nS_st7_b30_c1;
  assign nS_st8_b31_c1 = nS_st7_b31_c1;
  assign nS_st8_b32_c1 = nS_st7_b32_c1;
  assign nS_st8_b33_c1 = nS_st7_b33_c1;
  assign nS_st8_b34_c1 = nS_st7_b34_c1;
  assign nS_st8_b35_c1 = nS_st7_b35_c1;
  assign nS_st8_b36_c1 = nS_st7_b36_c1;
  assign nS_st8_b37_c1 = nS_st7_b37_c1;
  assign nS_st8_b38_c1 = nS_st7_b38_c1;
  assign nS_st8_b39_c1 = nS_st7_b39_c1;
  assign nS_st8_b40_c1 = nS_st7_b40_c1;
  assign nS_st8_b41_c1 = nS_st7_b41_c1;
  assign nS_st8_b42_c1 = nS_st7_b42_c1;
  assign nS_st8_b43_c1 = nS_st7_b43_c1;
  assign nS_st8_b44_c1 = nS_st7_b44_c1;
  assign nS_st8_b45_c1 = nS_st7_b45_c1;
  assign nS_st8_b46_c1 = nS_st7_b46_c1;
  assign nS_st8_b47_c1 = nS_st7_b47_c1;
  assign nS_st8_b48_c1 = nS_st7_b48_c1;
  assign nS_st8_b49_c1 = nS_st7_b49_c1;
  assign nS_st8_b50_c1 = nS_st7_b50_c1;
  assign nS_st8_b51_c1 = nS_st7_b51_c1;
  assign nS_st8_b52_c1 = nS_st7_b52_c1;
  assign nS_st8_b53_c1 = nS_st7_b53_c1;
  assign nS_st8_b54_c1 = nS_st7_b54_c1;
  assign nS_st8_b55_c1 = nS_st7_b55_c1;
  assign nS_st8_b56_c1 = nS_st7_b56_c1;
  assign nS_st8_b57_c1 = nS_st7_b57_c1;
  assign nS_st8_b58_c1 = nS_st7_b58_c1;
  assign nS_st8_b59_c1 = nS_st7_b59_c1;
  assign nS_st8_b60_c1 = nS_st7_b60_c1;
  assign nS_st8_b61_c1 = nS_st7_b61_c1;
  assign nS_st8_b62_c1 = nS_st7_b62_c1;
  assign nS_st8_b63_c1 = nS_st7_b63_c1;
  assign nS_st8_b64_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b64_c0 : nS_st7_b64_c1;
  assign nS_st8_b65_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b65_c0 : nS_st7_b65_c1;
  assign nS_st8_b66_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b66_c0 : nS_st7_b66_c1;
  assign nS_st8_b67_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b67_c0 : nS_st7_b67_c1;
  assign nS_st8_b68_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b68_c0 : nS_st7_b68_c1;
  assign nS_st8_b69_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b69_c0 : nS_st7_b69_c1;
  assign nS_st8_b70_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b70_c0 : nS_st7_b70_c1;
  assign nS_st8_b71_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b71_c0 : nS_st7_b71_c1;
  assign nS_st8_b72_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b72_c0 : nS_st7_b72_c1;
  assign nS_st8_b73_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b73_c0 : nS_st7_b73_c1;
  assign nS_st8_b74_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b74_c0 : nS_st7_b74_c1;
  assign nS_st8_b75_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b75_c0 : nS_st7_b75_c1;
  assign nS_st8_b76_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b76_c0 : nS_st7_b76_c1;
  assign nS_st8_b77_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b77_c0 : nS_st7_b77_c1;
  assign nS_st8_b78_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b78_c0 : nS_st7_b78_c1;
  assign nS_st8_b79_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b79_c0 : nS_st7_b79_c1;
  assign nS_st8_b80_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b80_c0 : nS_st7_b80_c1;
  assign nS_st8_b81_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b81_c0 : nS_st7_b81_c1;
  assign nS_st8_b82_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b82_c0 : nS_st7_b82_c1;
  assign nS_st8_b83_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b83_c0 : nS_st7_b83_c1;
  assign nS_st8_b84_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b84_c0 : nS_st7_b84_c1;
  assign nS_st8_b85_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b85_c0 : nS_st7_b85_c1;
  assign nS_st8_b86_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b86_c0 : nS_st7_b86_c1;
  assign nS_st8_b87_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b87_c0 : nS_st7_b87_c1;
  assign nS_st8_b88_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b88_c0 : nS_st7_b88_c1;
  assign nS_st8_b89_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b89_c0 : nS_st7_b89_c1;
  assign nS_st8_b90_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b90_c0 : nS_st7_b90_c1;
  assign nS_st8_b91_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b91_c0 : nS_st7_b91_c1;
  assign nS_st8_b92_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b92_c0 : nS_st7_b92_c1;
  assign nS_st8_b93_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b93_c0 : nS_st7_b93_c1;
  assign nS_st8_b94_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b94_c0 : nS_st7_b94_c1;
  assign nS_st8_b95_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b95_c0 : nS_st7_b95_c1;
  assign nS_st8_b96_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b96_c0 : nS_st7_b96_c1;
  assign nS_st8_b97_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b97_c0 : nS_st7_b97_c1;
  assign nS_st8_b98_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b98_c0 : nS_st7_b98_c1;
  assign nS_st8_b99_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b99_c0 : nS_st7_b99_c1;
  assign nS_st8_b100_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b100_c0 : nS_st7_b100_c1;
  assign nS_st8_b101_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b101_c0 : nS_st7_b101_c1;
  assign nS_st8_b102_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b102_c0 : nS_st7_b102_c1;
  assign nS_st8_b103_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b103_c0 : nS_st7_b103_c1;
  assign nS_st8_b104_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b104_c0 : nS_st7_b104_c1;
  assign nS_st8_b105_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b105_c0 : nS_st7_b105_c1;
  assign nS_st8_b106_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b106_c0 : nS_st7_b106_c1;
  assign nS_st8_b107_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b107_c0 : nS_st7_b107_c1;
  assign nS_st8_b108_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b108_c0 : nS_st7_b108_c1;
  assign nS_st8_b109_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b109_c0 : nS_st7_b109_c1;
  assign nS_st8_b110_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b110_c0 : nS_st7_b110_c1;
  assign nS_st8_b111_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b111_c0 : nS_st7_b111_c1;
  assign nS_st8_b112_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b112_c0 : nS_st7_b112_c1;
  assign nS_st8_b113_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b113_c0 : nS_st7_b113_c1;
  assign nS_st8_b114_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b114_c0 : nS_st7_b114_c1;
  assign nS_st8_b115_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b115_c0 : nS_st7_b115_c1;
  assign nS_st8_b116_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b116_c0 : nS_st7_b116_c1;
  assign nS_st8_b117_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b117_c0 : nS_st7_b117_c1;
  assign nS_st8_b118_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b118_c0 : nS_st7_b118_c1;
  assign nS_st8_b119_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b119_c0 : nS_st7_b119_c1;
  assign nS_st8_b120_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b120_c0 : nS_st7_b120_c1;
  assign nS_st8_b121_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b121_c0 : nS_st7_b121_c1;
  assign nS_st8_b122_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b122_c0 : nS_st7_b122_c1;
  assign nS_st8_b123_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b123_c0 : nS_st7_b123_c1;
  assign nS_st8_b124_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b124_c0 : nS_st7_b124_c1;
  assign nS_st8_b125_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b125_c0 : nS_st7_b125_c1;
  assign nS_st8_b126_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b126_c0 : nS_st7_b126_c1;
  assign nS_st8_b127_c1 = (nC_st7_b63_c1 == 0) ? nS_st7_b127_c0 : nS_st7_b127_c1;
  assign nC_st8_b127_c0 = (nC_st7_b63_c0 == 0) ? nC_st7_b127_c0 : nC_st7_b127_c1;
  assign nC_st8_b127_c1 = (nC_st7_b63_c1 == 0) ? nC_st7_b127_c0 : nC_st7_b127_c1;

  assign out_S[0] = (in_CI == 0) ? nS_st8_b0_c0 : nS_st8_b0_c1;
  assign out_S[1] = (in_CI == 0) ? nS_st8_b1_c0 : nS_st8_b1_c1;
  assign out_S[2] = (in_CI == 0) ? nS_st8_b2_c0 : nS_st8_b2_c1;
  assign out_S[3] = (in_CI == 0) ? nS_st8_b3_c0 : nS_st8_b3_c1;
  assign out_S[4] = (in_CI == 0) ? nS_st8_b4_c0 : nS_st8_b4_c1;
  assign out_S[5] = (in_CI == 0) ? nS_st8_b5_c0 : nS_st8_b5_c1;
  assign out_S[6] = (in_CI == 0) ? nS_st8_b6_c0 : nS_st8_b6_c1;
  assign out_S[7] = (in_CI == 0) ? nS_st8_b7_c0 : nS_st8_b7_c1;
  assign out_S[8] = (in_CI == 0) ? nS_st8_b8_c0 : nS_st8_b8_c1;
  assign out_S[9] = (in_CI == 0) ? nS_st8_b9_c0 : nS_st8_b9_c1;
  assign out_S[10] = (in_CI == 0) ? nS_st8_b10_c0 : nS_st8_b10_c1;
  assign out_S[11] = (in_CI == 0) ? nS_st8_b11_c0 : nS_st8_b11_c1;
  assign out_S[12] = (in_CI == 0) ? nS_st8_b12_c0 : nS_st8_b12_c1;
  assign out_S[13] = (in_CI == 0) ? nS_st8_b13_c0 : nS_st8_b13_c1;
  assign out_S[14] = (in_CI == 0) ? nS_st8_b14_c0 : nS_st8_b14_c1;
  assign out_S[15] = (in_CI == 0) ? nS_st8_b15_c0 : nS_st8_b15_c1;
  assign out_S[16] = (in_CI == 0) ? nS_st8_b16_c0 : nS_st8_b16_c1;
  assign out_S[17] = (in_CI == 0) ? nS_st8_b17_c0 : nS_st8_b17_c1;
  assign out_S[18] = (in_CI == 0) ? nS_st8_b18_c0 : nS_st8_b18_c1;
  assign out_S[19] = (in_CI == 0) ? nS_st8_b19_c0 : nS_st8_b19_c1;
  assign out_S[20] = (in_CI == 0) ? nS_st8_b20_c0 : nS_st8_b20_c1;
  assign out_S[21] = (in_CI == 0) ? nS_st8_b21_c0 : nS_st8_b21_c1;
  assign out_S[22] = (in_CI == 0) ? nS_st8_b22_c0 : nS_st8_b22_c1;
  assign out_S[23] = (in_CI == 0) ? nS_st8_b23_c0 : nS_st8_b23_c1;
  assign out_S[24] = (in_CI == 0) ? nS_st8_b24_c0 : nS_st8_b24_c1;
  assign out_S[25] = (in_CI == 0) ? nS_st8_b25_c0 : nS_st8_b25_c1;
  assign out_S[26] = (in_CI == 0) ? nS_st8_b26_c0 : nS_st8_b26_c1;
  assign out_S[27] = (in_CI == 0) ? nS_st8_b27_c0 : nS_st8_b27_c1;
  assign out_S[28] = (in_CI == 0) ? nS_st8_b28_c0 : nS_st8_b28_c1;
  assign out_S[29] = (in_CI == 0) ? nS_st8_b29_c0 : nS_st8_b29_c1;
  assign out_S[30] = (in_CI == 0) ? nS_st8_b30_c0 : nS_st8_b30_c1;
  assign out_S[31] = (in_CI == 0) ? nS_st8_b31_c0 : nS_st8_b31_c1;
  assign out_S[32] = (in_CI == 0) ? nS_st8_b32_c0 : nS_st8_b32_c1;
  assign out_S[33] = (in_CI == 0) ? nS_st8_b33_c0 : nS_st8_b33_c1;
  assign out_S[34] = (in_CI == 0) ? nS_st8_b34_c0 : nS_st8_b34_c1;
  assign out_S[35] = (in_CI == 0) ? nS_st8_b35_c0 : nS_st8_b35_c1;
  assign out_S[36] = (in_CI == 0) ? nS_st8_b36_c0 : nS_st8_b36_c1;
  assign out_S[37] = (in_CI == 0) ? nS_st8_b37_c0 : nS_st8_b37_c1;
  assign out_S[38] = (in_CI == 0) ? nS_st8_b38_c0 : nS_st8_b38_c1;
  assign out_S[39] = (in_CI == 0) ? nS_st8_b39_c0 : nS_st8_b39_c1;
  assign out_S[40] = (in_CI == 0) ? nS_st8_b40_c0 : nS_st8_b40_c1;
  assign out_S[41] = (in_CI == 0) ? nS_st8_b41_c0 : nS_st8_b41_c1;
  assign out_S[42] = (in_CI == 0) ? nS_st8_b42_c0 : nS_st8_b42_c1;
  assign out_S[43] = (in_CI == 0) ? nS_st8_b43_c0 : nS_st8_b43_c1;
  assign out_S[44] = (in_CI == 0) ? nS_st8_b44_c0 : nS_st8_b44_c1;
  assign out_S[45] = (in_CI == 0) ? nS_st8_b45_c0 : nS_st8_b45_c1;
  assign out_S[46] = (in_CI == 0) ? nS_st8_b46_c0 : nS_st8_b46_c1;
  assign out_S[47] = (in_CI == 0) ? nS_st8_b47_c0 : nS_st8_b47_c1;
  assign out_S[48] = (in_CI == 0) ? nS_st8_b48_c0 : nS_st8_b48_c1;
  assign out_S[49] = (in_CI == 0) ? nS_st8_b49_c0 : nS_st8_b49_c1;
  assign out_S[50] = (in_CI == 0) ? nS_st8_b50_c0 : nS_st8_b50_c1;
  assign out_S[51] = (in_CI == 0) ? nS_st8_b51_c0 : nS_st8_b51_c1;
  assign out_S[52] = (in_CI == 0) ? nS_st8_b52_c0 : nS_st8_b52_c1;
  assign out_S[53] = (in_CI == 0) ? nS_st8_b53_c0 : nS_st8_b53_c1;
  assign out_S[54] = (in_CI == 0) ? nS_st8_b54_c0 : nS_st8_b54_c1;
  assign out_S[55] = (in_CI == 0) ? nS_st8_b55_c0 : nS_st8_b55_c1;
  assign out_S[56] = (in_CI == 0) ? nS_st8_b56_c0 : nS_st8_b56_c1;
  assign out_S[57] = (in_CI == 0) ? nS_st8_b57_c0 : nS_st8_b57_c1;
  assign out_S[58] = (in_CI == 0) ? nS_st8_b58_c0 : nS_st8_b58_c1;
  assign out_S[59] = (in_CI == 0) ? nS_st8_b59_c0 : nS_st8_b59_c1;
  assign out_S[60] = (in_CI == 0) ? nS_st8_b60_c0 : nS_st8_b60_c1;
  assign out_S[61] = (in_CI == 0) ? nS_st8_b61_c0 : nS_st8_b61_c1;
  assign out_S[62] = (in_CI == 0) ? nS_st8_b62_c0 : nS_st8_b62_c1;
  assign out_S[63] = (in_CI == 0) ? nS_st8_b63_c0 : nS_st8_b63_c1;
  assign out_S[64] = (in_CI == 0) ? nS_st8_b64_c0 : nS_st8_b64_c1;
  assign out_S[65] = (in_CI == 0) ? nS_st8_b65_c0 : nS_st8_b65_c1;
  assign out_S[66] = (in_CI == 0) ? nS_st8_b66_c0 : nS_st8_b66_c1;
  assign out_S[67] = (in_CI == 0) ? nS_st8_b67_c0 : nS_st8_b67_c1;
  assign out_S[68] = (in_CI == 0) ? nS_st8_b68_c0 : nS_st8_b68_c1;
  assign out_S[69] = (in_CI == 0) ? nS_st8_b69_c0 : nS_st8_b69_c1;
  assign out_S[70] = (in_CI == 0) ? nS_st8_b70_c0 : nS_st8_b70_c1;
  assign out_S[71] = (in_CI == 0) ? nS_st8_b71_c0 : nS_st8_b71_c1;
  assign out_S[72] = (in_CI == 0) ? nS_st8_b72_c0 : nS_st8_b72_c1;
  assign out_S[73] = (in_CI == 0) ? nS_st8_b73_c0 : nS_st8_b73_c1;
  assign out_S[74] = (in_CI == 0) ? nS_st8_b74_c0 : nS_st8_b74_c1;
  assign out_S[75] = (in_CI == 0) ? nS_st8_b75_c0 : nS_st8_b75_c1;
  assign out_S[76] = (in_CI == 0) ? nS_st8_b76_c0 : nS_st8_b76_c1;
  assign out_S[77] = (in_CI == 0) ? nS_st8_b77_c0 : nS_st8_b77_c1;
  assign out_S[78] = (in_CI == 0) ? nS_st8_b78_c0 : nS_st8_b78_c1;
  assign out_S[79] = (in_CI == 0) ? nS_st8_b79_c0 : nS_st8_b79_c1;
  assign out_S[80] = (in_CI == 0) ? nS_st8_b80_c0 : nS_st8_b80_c1;
  assign out_S[81] = (in_CI == 0) ? nS_st8_b81_c0 : nS_st8_b81_c1;
  assign out_S[82] = (in_CI == 0) ? nS_st8_b82_c0 : nS_st8_b82_c1;
  assign out_S[83] = (in_CI == 0) ? nS_st8_b83_c0 : nS_st8_b83_c1;
  assign out_S[84] = (in_CI == 0) ? nS_st8_b84_c0 : nS_st8_b84_c1;
  assign out_S[85] = (in_CI == 0) ? nS_st8_b85_c0 : nS_st8_b85_c1;
  assign out_S[86] = (in_CI == 0) ? nS_st8_b86_c0 : nS_st8_b86_c1;
  assign out_S[87] = (in_CI == 0) ? nS_st8_b87_c0 : nS_st8_b87_c1;
  assign out_S[88] = (in_CI == 0) ? nS_st8_b88_c0 : nS_st8_b88_c1;
  assign out_S[89] = (in_CI == 0) ? nS_st8_b89_c0 : nS_st8_b89_c1;
  assign out_S[90] = (in_CI == 0) ? nS_st8_b90_c0 : nS_st8_b90_c1;
  assign out_S[91] = (in_CI == 0) ? nS_st8_b91_c0 : nS_st8_b91_c1;
  assign out_S[92] = (in_CI == 0) ? nS_st8_b92_c0 : nS_st8_b92_c1;
  assign out_S[93] = (in_CI == 0) ? nS_st8_b93_c0 : nS_st8_b93_c1;
  assign out_S[94] = (in_CI == 0) ? nS_st8_b94_c0 : nS_st8_b94_c1;
  assign out_S[95] = (in_CI == 0) ? nS_st8_b95_c0 : nS_st8_b95_c1;
  assign out_S[96] = (in_CI == 0) ? nS_st8_b96_c0 : nS_st8_b96_c1;
  assign out_S[97] = (in_CI == 0) ? nS_st8_b97_c0 : nS_st8_b97_c1;
  assign out_S[98] = (in_CI == 0) ? nS_st8_b98_c0 : nS_st8_b98_c1;
  assign out_S[99] = (in_CI == 0) ? nS_st8_b99_c0 : nS_st8_b99_c1;
  assign out_S[100] = (in_CI == 0) ? nS_st8_b100_c0 : nS_st8_b100_c1;
  assign out_S[101] = (in_CI == 0) ? nS_st8_b101_c0 : nS_st8_b101_c1;
  assign out_S[102] = (in_CI == 0) ? nS_st8_b102_c0 : nS_st8_b102_c1;
  assign out_S[103] = (in_CI == 0) ? nS_st8_b103_c0 : nS_st8_b103_c1;
  assign out_S[104] = (in_CI == 0) ? nS_st8_b104_c0 : nS_st8_b104_c1;
  assign out_S[105] = (in_CI == 0) ? nS_st8_b105_c0 : nS_st8_b105_c1;
  assign out_S[106] = (in_CI == 0) ? nS_st8_b106_c0 : nS_st8_b106_c1;
  assign out_S[107] = (in_CI == 0) ? nS_st8_b107_c0 : nS_st8_b107_c1;
  assign out_S[108] = (in_CI == 0) ? nS_st8_b108_c0 : nS_st8_b108_c1;
  assign out_S[109] = (in_CI == 0) ? nS_st8_b109_c0 : nS_st8_b109_c1;
  assign out_S[110] = (in_CI == 0) ? nS_st8_b110_c0 : nS_st8_b110_c1;
  assign out_S[111] = (in_CI == 0) ? nS_st8_b111_c0 : nS_st8_b111_c1;
  assign out_S[112] = (in_CI == 0) ? nS_st8_b112_c0 : nS_st8_b112_c1;
  assign out_S[113] = (in_CI == 0) ? nS_st8_b113_c0 : nS_st8_b113_c1;
  assign out_S[114] = (in_CI == 0) ? nS_st8_b114_c0 : nS_st8_b114_c1;
  assign out_S[115] = (in_CI == 0) ? nS_st8_b115_c0 : nS_st8_b115_c1;
  assign out_S[116] = (in_CI == 0) ? nS_st8_b116_c0 : nS_st8_b116_c1;
  assign out_S[117] = (in_CI == 0) ? nS_st8_b117_c0 : nS_st8_b117_c1;
  assign out_S[118] = (in_CI == 0) ? nS_st8_b118_c0 : nS_st8_b118_c1;
  assign out_S[119] = (in_CI == 0) ? nS_st8_b119_c0 : nS_st8_b119_c1;
  assign out_S[120] = (in_CI == 0) ? nS_st8_b120_c0 : nS_st8_b120_c1;
  assign out_S[121] = (in_CI == 0) ? nS_st8_b121_c0 : nS_st8_b121_c1;
  assign out_S[122] = (in_CI == 0) ? nS_st8_b122_c0 : nS_st8_b122_c1;
  assign out_S[123] = (in_CI == 0) ? nS_st8_b123_c0 : nS_st8_b123_c1;
  assign out_S[124] = (in_CI == 0) ? nS_st8_b124_c0 : nS_st8_b124_c1;
  assign out_S[125] = (in_CI == 0) ? nS_st8_b125_c0 : nS_st8_b125_c1;
  assign out_S[126] = (in_CI == 0) ? nS_st8_b126_c0 : nS_st8_b126_c1;
  assign out_S[127] = (in_CI == 0) ? nS_st8_b127_c0 : nS_st8_b127_c1;
  assign out_CO = (in_CI == 0) ? nC_st8_b127_c0 : nC_st8_b127_c1;
endmodule

