module VKSA_64 (in_A, in_B, in_CI, out_S, out_CO);
  input [63:0] in_A, in_B;
  input in_CI;
  output [63:0] out_S;
  output out_CO;

  assign nG_0_0 = in_A[0] & in_B[0];
  assign nP_0_0 = in_A[0] ^ in_B[0];
  assign nG_1_1 = in_A[1] & in_B[1];
  assign nP_1_1 = in_A[1] ^ in_B[1];
  assign nG_2_2 = in_A[2] & in_B[2];
  assign nP_2_2 = in_A[2] ^ in_B[2];
  assign nG_3_3 = in_A[3] & in_B[3];
  assign nP_3_3 = in_A[3] ^ in_B[3];
  assign nG_4_4 = in_A[4] & in_B[4];
  assign nP_4_4 = in_A[4] ^ in_B[4];
  assign nG_5_5 = in_A[5] & in_B[5];
  assign nP_5_5 = in_A[5] ^ in_B[5];
  assign nG_6_6 = in_A[6] & in_B[6];
  assign nP_6_6 = in_A[6] ^ in_B[6];
  assign nG_7_7 = in_A[7] & in_B[7];
  assign nP_7_7 = in_A[7] ^ in_B[7];
  assign nG_8_8 = in_A[8] & in_B[8];
  assign nP_8_8 = in_A[8] ^ in_B[8];
  assign nG_9_9 = in_A[9] & in_B[9];
  assign nP_9_9 = in_A[9] ^ in_B[9];
  assign nG_10_10 = in_A[10] & in_B[10];
  assign nP_10_10 = in_A[10] ^ in_B[10];
  assign nG_11_11 = in_A[11] & in_B[11];
  assign nP_11_11 = in_A[11] ^ in_B[11];
  assign nG_12_12 = in_A[12] & in_B[12];
  assign nP_12_12 = in_A[12] ^ in_B[12];
  assign nG_13_13 = in_A[13] & in_B[13];
  assign nP_13_13 = in_A[13] ^ in_B[13];
  assign nG_14_14 = in_A[14] & in_B[14];
  assign nP_14_14 = in_A[14] ^ in_B[14];
  assign nG_15_15 = in_A[15] & in_B[15];
  assign nP_15_15 = in_A[15] ^ in_B[15];
  assign nG_16_16 = in_A[16] & in_B[16];
  assign nP_16_16 = in_A[16] ^ in_B[16];
  assign nG_17_17 = in_A[17] & in_B[17];
  assign nP_17_17 = in_A[17] ^ in_B[17];
  assign nG_18_18 = in_A[18] & in_B[18];
  assign nP_18_18 = in_A[18] ^ in_B[18];
  assign nG_19_19 = in_A[19] & in_B[19];
  assign nP_19_19 = in_A[19] ^ in_B[19];
  assign nG_20_20 = in_A[20] & in_B[20];
  assign nP_20_20 = in_A[20] ^ in_B[20];
  assign nG_21_21 = in_A[21] & in_B[21];
  assign nP_21_21 = in_A[21] ^ in_B[21];
  assign nG_22_22 = in_A[22] & in_B[22];
  assign nP_22_22 = in_A[22] ^ in_B[22];
  assign nG_23_23 = in_A[23] & in_B[23];
  assign nP_23_23 = in_A[23] ^ in_B[23];
  assign nG_24_24 = in_A[24] & in_B[24];
  assign nP_24_24 = in_A[24] ^ in_B[24];
  assign nG_25_25 = in_A[25] & in_B[25];
  assign nP_25_25 = in_A[25] ^ in_B[25];
  assign nG_26_26 = in_A[26] & in_B[26];
  assign nP_26_26 = in_A[26] ^ in_B[26];
  assign nG_27_27 = in_A[27] & in_B[27];
  assign nP_27_27 = in_A[27] ^ in_B[27];
  assign nG_28_28 = in_A[28] & in_B[28];
  assign nP_28_28 = in_A[28] ^ in_B[28];
  assign nG_29_29 = in_A[29] & in_B[29];
  assign nP_29_29 = in_A[29] ^ in_B[29];
  assign nG_30_30 = in_A[30] & in_B[30];
  assign nP_30_30 = in_A[30] ^ in_B[30];
  assign nG_31_31 = in_A[31] & in_B[31];
  assign nP_31_31 = in_A[31] ^ in_B[31];
  assign nG_32_32 = in_A[32] & in_B[32];
  assign nP_32_32 = in_A[32] ^ in_B[32];
  assign nG_33_33 = in_A[33] & in_B[33];
  assign nP_33_33 = in_A[33] ^ in_B[33];
  assign nG_34_34 = in_A[34] & in_B[34];
  assign nP_34_34 = in_A[34] ^ in_B[34];
  assign nG_35_35 = in_A[35] & in_B[35];
  assign nP_35_35 = in_A[35] ^ in_B[35];
  assign nG_36_36 = in_A[36] & in_B[36];
  assign nP_36_36 = in_A[36] ^ in_B[36];
  assign nG_37_37 = in_A[37] & in_B[37];
  assign nP_37_37 = in_A[37] ^ in_B[37];
  assign nG_38_38 = in_A[38] & in_B[38];
  assign nP_38_38 = in_A[38] ^ in_B[38];
  assign nG_39_39 = in_A[39] & in_B[39];
  assign nP_39_39 = in_A[39] ^ in_B[39];
  assign nG_40_40 = in_A[40] & in_B[40];
  assign nP_40_40 = in_A[40] ^ in_B[40];
  assign nG_41_41 = in_A[41] & in_B[41];
  assign nP_41_41 = in_A[41] ^ in_B[41];
  assign nG_42_42 = in_A[42] & in_B[42];
  assign nP_42_42 = in_A[42] ^ in_B[42];
  assign nG_43_43 = in_A[43] & in_B[43];
  assign nP_43_43 = in_A[43] ^ in_B[43];
  assign nG_44_44 = in_A[44] & in_B[44];
  assign nP_44_44 = in_A[44] ^ in_B[44];
  assign nG_45_45 = in_A[45] & in_B[45];
  assign nP_45_45 = in_A[45] ^ in_B[45];
  assign nG_46_46 = in_A[46] & in_B[46];
  assign nP_46_46 = in_A[46] ^ in_B[46];
  assign nG_47_47 = in_A[47] & in_B[47];
  assign nP_47_47 = in_A[47] ^ in_B[47];
  assign nG_48_48 = in_A[48] & in_B[48];
  assign nP_48_48 = in_A[48] ^ in_B[48];
  assign nG_49_49 = in_A[49] & in_B[49];
  assign nP_49_49 = in_A[49] ^ in_B[49];
  assign nG_50_50 = in_A[50] & in_B[50];
  assign nP_50_50 = in_A[50] ^ in_B[50];
  assign nG_51_51 = in_A[51] & in_B[51];
  assign nP_51_51 = in_A[51] ^ in_B[51];
  assign nG_52_52 = in_A[52] & in_B[52];
  assign nP_52_52 = in_A[52] ^ in_B[52];
  assign nG_53_53 = in_A[53] & in_B[53];
  assign nP_53_53 = in_A[53] ^ in_B[53];
  assign nG_54_54 = in_A[54] & in_B[54];
  assign nP_54_54 = in_A[54] ^ in_B[54];
  assign nG_55_55 = in_A[55] & in_B[55];
  assign nP_55_55 = in_A[55] ^ in_B[55];
  assign nG_56_56 = in_A[56] & in_B[56];
  assign nP_56_56 = in_A[56] ^ in_B[56];
  assign nG_57_57 = in_A[57] & in_B[57];
  assign nP_57_57 = in_A[57] ^ in_B[57];
  assign nG_58_58 = in_A[58] & in_B[58];
  assign nP_58_58 = in_A[58] ^ in_B[58];
  assign nG_59_59 = in_A[59] & in_B[59];
  assign nP_59_59 = in_A[59] ^ in_B[59];
  assign nG_60_60 = in_A[60] & in_B[60];
  assign nP_60_60 = in_A[60] ^ in_B[60];
  assign nG_61_61 = in_A[61] & in_B[61];
  assign nP_61_61 = in_A[61] ^ in_B[61];
  assign nG_62_62 = in_A[62] & in_B[62];
  assign nP_62_62 = in_A[62] ^ in_B[62];
  assign nG_63_63 = in_A[63] & in_B[63];
  assign nP_63_63 = in_A[63] ^ in_B[63];

  assign nG_63_62 = nG_63_63 | (nP_63_63 & nG_62_62);
  assign nP_63_62 = nP_63_63 & nP_62_62;
  assign nG_62_61 = nG_62_62 | (nP_62_62 & nG_61_61);
  assign nP_62_61 = nP_62_62 & nP_61_61;
  assign nG_61_60 = nG_61_61 | (nP_61_61 & nG_60_60);
  assign nP_61_60 = nP_61_61 & nP_60_60;
  assign nG_60_59 = nG_60_60 | (nP_60_60 & nG_59_59);
  assign nP_60_59 = nP_60_60 & nP_59_59;
  assign nG_59_58 = nG_59_59 | (nP_59_59 & nG_58_58);
  assign nP_59_58 = nP_59_59 & nP_58_58;
  assign nG_58_57 = nG_58_58 | (nP_58_58 & nG_57_57);
  assign nP_58_57 = nP_58_58 & nP_57_57;
  assign nG_57_56 = nG_57_57 | (nP_57_57 & nG_56_56);
  assign nP_57_56 = nP_57_57 & nP_56_56;
  assign nG_56_55 = nG_56_56 | (nP_56_56 & nG_55_55);
  assign nP_56_55 = nP_56_56 & nP_55_55;
  assign nG_55_54 = nG_55_55 | (nP_55_55 & nG_54_54);
  assign nP_55_54 = nP_55_55 & nP_54_54;
  assign nG_54_53 = nG_54_54 | (nP_54_54 & nG_53_53);
  assign nP_54_53 = nP_54_54 & nP_53_53;
  assign nG_53_52 = nG_53_53 | (nP_53_53 & nG_52_52);
  assign nP_53_52 = nP_53_53 & nP_52_52;
  assign nG_52_51 = nG_52_52 | (nP_52_52 & nG_51_51);
  assign nP_52_51 = nP_52_52 & nP_51_51;
  assign nG_51_50 = nG_51_51 | (nP_51_51 & nG_50_50);
  assign nP_51_50 = nP_51_51 & nP_50_50;
  assign nG_50_49 = nG_50_50 | (nP_50_50 & nG_49_49);
  assign nP_50_49 = nP_50_50 & nP_49_49;
  assign nG_49_48 = nG_49_49 | (nP_49_49 & nG_48_48);
  assign nP_49_48 = nP_49_49 & nP_48_48;
  assign nG_48_47 = nG_48_48 | (nP_48_48 & nG_47_47);
  assign nP_48_47 = nP_48_48 & nP_47_47;
  assign nG_47_46 = nG_47_47 | (nP_47_47 & nG_46_46);
  assign nP_47_46 = nP_47_47 & nP_46_46;
  assign nG_46_45 = nG_46_46 | (nP_46_46 & nG_45_45);
  assign nP_46_45 = nP_46_46 & nP_45_45;
  assign nG_45_44 = nG_45_45 | (nP_45_45 & nG_44_44);
  assign nP_45_44 = nP_45_45 & nP_44_44;
  assign nG_44_43 = nG_44_44 | (nP_44_44 & nG_43_43);
  assign nP_44_43 = nP_44_44 & nP_43_43;
  assign nG_43_42 = nG_43_43 | (nP_43_43 & nG_42_42);
  assign nP_43_42 = nP_43_43 & nP_42_42;
  assign nG_42_41 = nG_42_42 | (nP_42_42 & nG_41_41);
  assign nP_42_41 = nP_42_42 & nP_41_41;
  assign nG_41_40 = nG_41_41 | (nP_41_41 & nG_40_40);
  assign nP_41_40 = nP_41_41 & nP_40_40;
  assign nG_40_39 = nG_40_40 | (nP_40_40 & nG_39_39);
  assign nP_40_39 = nP_40_40 & nP_39_39;
  assign nG_39_38 = nG_39_39 | (nP_39_39 & nG_38_38);
  assign nP_39_38 = nP_39_39 & nP_38_38;
  assign nG_38_37 = nG_38_38 | (nP_38_38 & nG_37_37);
  assign nP_38_37 = nP_38_38 & nP_37_37;
  assign nG_37_36 = nG_37_37 | (nP_37_37 & nG_36_36);
  assign nP_37_36 = nP_37_37 & nP_36_36;
  assign nG_36_35 = nG_36_36 | (nP_36_36 & nG_35_35);
  assign nP_36_35 = nP_36_36 & nP_35_35;
  assign nG_35_34 = nG_35_35 | (nP_35_35 & nG_34_34);
  assign nP_35_34 = nP_35_35 & nP_34_34;
  assign nG_34_33 = nG_34_34 | (nP_34_34 & nG_33_33);
  assign nP_34_33 = nP_34_34 & nP_33_33;
  assign nG_33_32 = nG_33_33 | (nP_33_33 & nG_32_32);
  assign nP_33_32 = nP_33_33 & nP_32_32;
  assign nG_32_31 = nG_32_32 | (nP_32_32 & nG_31_31);
  assign nP_32_31 = nP_32_32 & nP_31_31;
  assign nG_31_30 = nG_31_31 | (nP_31_31 & nG_30_30);
  assign nP_31_30 = nP_31_31 & nP_30_30;
  assign nG_30_29 = nG_30_30 | (nP_30_30 & nG_29_29);
  assign nP_30_29 = nP_30_30 & nP_29_29;
  assign nG_29_28 = nG_29_29 | (nP_29_29 & nG_28_28);
  assign nP_29_28 = nP_29_29 & nP_28_28;
  assign nG_28_27 = nG_28_28 | (nP_28_28 & nG_27_27);
  assign nP_28_27 = nP_28_28 & nP_27_27;
  assign nG_27_26 = nG_27_27 | (nP_27_27 & nG_26_26);
  assign nP_27_26 = nP_27_27 & nP_26_26;
  assign nG_26_25 = nG_26_26 | (nP_26_26 & nG_25_25);
  assign nP_26_25 = nP_26_26 & nP_25_25;
  assign nG_25_24 = nG_25_25 | (nP_25_25 & nG_24_24);
  assign nP_25_24 = nP_25_25 & nP_24_24;
  assign nG_24_23 = nG_24_24 | (nP_24_24 & nG_23_23);
  assign nP_24_23 = nP_24_24 & nP_23_23;
  assign nG_23_22 = nG_23_23 | (nP_23_23 & nG_22_22);
  assign nP_23_22 = nP_23_23 & nP_22_22;
  assign nG_22_21 = nG_22_22 | (nP_22_22 & nG_21_21);
  assign nP_22_21 = nP_22_22 & nP_21_21;
  assign nG_21_20 = nG_21_21 | (nP_21_21 & nG_20_20);
  assign nP_21_20 = nP_21_21 & nP_20_20;
  assign nG_20_19 = nG_20_20 | (nP_20_20 & nG_19_19);
  assign nP_20_19 = nP_20_20 & nP_19_19;
  assign nG_19_18 = nG_19_19 | (nP_19_19 & nG_18_18);
  assign nP_19_18 = nP_19_19 & nP_18_18;
  assign nG_18_17 = nG_18_18 | (nP_18_18 & nG_17_17);
  assign nP_18_17 = nP_18_18 & nP_17_17;
  assign nG_17_16 = nG_17_17 | (nP_17_17 & nG_16_16);
  assign nP_17_16 = nP_17_17 & nP_16_16;
  assign nG_16_15 = nG_16_16 | (nP_16_16 & nG_15_15);
  assign nP_16_15 = nP_16_16 & nP_15_15;
  assign nG_15_14 = nG_15_15 | (nP_15_15 & nG_14_14);
  assign nP_15_14 = nP_15_15 & nP_14_14;
  assign nG_14_13 = nG_14_14 | (nP_14_14 & nG_13_13);
  assign nP_14_13 = nP_14_14 & nP_13_13;
  assign nG_13_12 = nG_13_13 | (nP_13_13 & nG_12_12);
  assign nP_13_12 = nP_13_13 & nP_12_12;
  assign nG_12_11 = nG_12_12 | (nP_12_12 & nG_11_11);
  assign nP_12_11 = nP_12_12 & nP_11_11;
  assign nG_11_10 = nG_11_11 | (nP_11_11 & nG_10_10);
  assign nP_11_10 = nP_11_11 & nP_10_10;
  assign nG_10_9 = nG_10_10 | (nP_10_10 & nG_9_9);
  assign nP_10_9 = nP_10_10 & nP_9_9;
  assign nG_9_8 = nG_9_9 | (nP_9_9 & nG_8_8);
  assign nP_9_8 = nP_9_9 & nP_8_8;
  assign nG_8_7 = nG_8_8 | (nP_8_8 & nG_7_7);
  assign nP_8_7 = nP_8_8 & nP_7_7;
  assign nG_7_6 = nG_7_7 | (nP_7_7 & nG_6_6);
  assign nP_7_6 = nP_7_7 & nP_6_6;
  assign nG_6_5 = nG_6_6 | (nP_6_6 & nG_5_5);
  assign nP_6_5 = nP_6_6 & nP_5_5;
  assign nG_5_4 = nG_5_5 | (nP_5_5 & nG_4_4);
  assign nP_5_4 = nP_5_5 & nP_4_4;
  assign nG_4_3 = nG_4_4 | (nP_4_4 & nG_3_3);
  assign nP_4_3 = nP_4_4 & nP_3_3;
  assign nG_3_2 = nG_3_3 | (nP_3_3 & nG_2_2);
  assign nP_3_2 = nP_3_3 & nP_2_2;
  assign nG_2_1 = nG_2_2 | (nP_2_2 & nG_1_1);
  assign nP_2_1 = nP_2_2 & nP_1_1;
  assign nG_1_0 = nG_1_1 | (nP_1_1 & nG_0_0);
  assign nP_1_0 = nP_1_1 & nP_0_0;

  assign nG_63_60 = nG_63_62 | (nP_63_62 & nG_61_60);
  assign nP_63_60 = nP_63_62 & nP_61_60;
  assign nG_62_59 = nG_62_61 | (nP_62_61 & nG_60_59);
  assign nP_62_59 = nP_62_61 & nP_60_59;
  assign nG_61_58 = nG_61_60 | (nP_61_60 & nG_59_58);
  assign nP_61_58 = nP_61_60 & nP_59_58;
  assign nG_60_57 = nG_60_59 | (nP_60_59 & nG_58_57);
  assign nP_60_57 = nP_60_59 & nP_58_57;
  assign nG_59_56 = nG_59_58 | (nP_59_58 & nG_57_56);
  assign nP_59_56 = nP_59_58 & nP_57_56;
  assign nG_58_55 = nG_58_57 | (nP_58_57 & nG_56_55);
  assign nP_58_55 = nP_58_57 & nP_56_55;
  assign nG_57_54 = nG_57_56 | (nP_57_56 & nG_55_54);
  assign nP_57_54 = nP_57_56 & nP_55_54;
  assign nG_56_53 = nG_56_55 | (nP_56_55 & nG_54_53);
  assign nP_56_53 = nP_56_55 & nP_54_53;
  assign nG_55_52 = nG_55_54 | (nP_55_54 & nG_53_52);
  assign nP_55_52 = nP_55_54 & nP_53_52;
  assign nG_54_51 = nG_54_53 | (nP_54_53 & nG_52_51);
  assign nP_54_51 = nP_54_53 & nP_52_51;
  assign nG_53_50 = nG_53_52 | (nP_53_52 & nG_51_50);
  assign nP_53_50 = nP_53_52 & nP_51_50;
  assign nG_52_49 = nG_52_51 | (nP_52_51 & nG_50_49);
  assign nP_52_49 = nP_52_51 & nP_50_49;
  assign nG_51_48 = nG_51_50 | (nP_51_50 & nG_49_48);
  assign nP_51_48 = nP_51_50 & nP_49_48;
  assign nG_50_47 = nG_50_49 | (nP_50_49 & nG_48_47);
  assign nP_50_47 = nP_50_49 & nP_48_47;
  assign nG_49_46 = nG_49_48 | (nP_49_48 & nG_47_46);
  assign nP_49_46 = nP_49_48 & nP_47_46;
  assign nG_48_45 = nG_48_47 | (nP_48_47 & nG_46_45);
  assign nP_48_45 = nP_48_47 & nP_46_45;
  assign nG_47_44 = nG_47_46 | (nP_47_46 & nG_45_44);
  assign nP_47_44 = nP_47_46 & nP_45_44;
  assign nG_46_43 = nG_46_45 | (nP_46_45 & nG_44_43);
  assign nP_46_43 = nP_46_45 & nP_44_43;
  assign nG_45_42 = nG_45_44 | (nP_45_44 & nG_43_42);
  assign nP_45_42 = nP_45_44 & nP_43_42;
  assign nG_44_41 = nG_44_43 | (nP_44_43 & nG_42_41);
  assign nP_44_41 = nP_44_43 & nP_42_41;
  assign nG_43_40 = nG_43_42 | (nP_43_42 & nG_41_40);
  assign nP_43_40 = nP_43_42 & nP_41_40;
  assign nG_42_39 = nG_42_41 | (nP_42_41 & nG_40_39);
  assign nP_42_39 = nP_42_41 & nP_40_39;
  assign nG_41_38 = nG_41_40 | (nP_41_40 & nG_39_38);
  assign nP_41_38 = nP_41_40 & nP_39_38;
  assign nG_40_37 = nG_40_39 | (nP_40_39 & nG_38_37);
  assign nP_40_37 = nP_40_39 & nP_38_37;
  assign nG_39_36 = nG_39_38 | (nP_39_38 & nG_37_36);
  assign nP_39_36 = nP_39_38 & nP_37_36;
  assign nG_38_35 = nG_38_37 | (nP_38_37 & nG_36_35);
  assign nP_38_35 = nP_38_37 & nP_36_35;
  assign nG_37_34 = nG_37_36 | (nP_37_36 & nG_35_34);
  assign nP_37_34 = nP_37_36 & nP_35_34;
  assign nG_36_33 = nG_36_35 | (nP_36_35 & nG_34_33);
  assign nP_36_33 = nP_36_35 & nP_34_33;
  assign nG_35_32 = nG_35_34 | (nP_35_34 & nG_33_32);
  assign nP_35_32 = nP_35_34 & nP_33_32;
  assign nG_34_31 = nG_34_33 | (nP_34_33 & nG_32_31);
  assign nP_34_31 = nP_34_33 & nP_32_31;
  assign nG_33_30 = nG_33_32 | (nP_33_32 & nG_31_30);
  assign nP_33_30 = nP_33_32 & nP_31_30;
  assign nG_32_29 = nG_32_31 | (nP_32_31 & nG_30_29);
  assign nP_32_29 = nP_32_31 & nP_30_29;
  assign nG_31_28 = nG_31_30 | (nP_31_30 & nG_29_28);
  assign nP_31_28 = nP_31_30 & nP_29_28;
  assign nG_30_27 = nG_30_29 | (nP_30_29 & nG_28_27);
  assign nP_30_27 = nP_30_29 & nP_28_27;
  assign nG_29_26 = nG_29_28 | (nP_29_28 & nG_27_26);
  assign nP_29_26 = nP_29_28 & nP_27_26;
  assign nG_28_25 = nG_28_27 | (nP_28_27 & nG_26_25);
  assign nP_28_25 = nP_28_27 & nP_26_25;
  assign nG_27_24 = nG_27_26 | (nP_27_26 & nG_25_24);
  assign nP_27_24 = nP_27_26 & nP_25_24;
  assign nG_26_23 = nG_26_25 | (nP_26_25 & nG_24_23);
  assign nP_26_23 = nP_26_25 & nP_24_23;
  assign nG_25_22 = nG_25_24 | (nP_25_24 & nG_23_22);
  assign nP_25_22 = nP_25_24 & nP_23_22;
  assign nG_24_21 = nG_24_23 | (nP_24_23 & nG_22_21);
  assign nP_24_21 = nP_24_23 & nP_22_21;
  assign nG_23_20 = nG_23_22 | (nP_23_22 & nG_21_20);
  assign nP_23_20 = nP_23_22 & nP_21_20;
  assign nG_22_19 = nG_22_21 | (nP_22_21 & nG_20_19);
  assign nP_22_19 = nP_22_21 & nP_20_19;
  assign nG_21_18 = nG_21_20 | (nP_21_20 & nG_19_18);
  assign nP_21_18 = nP_21_20 & nP_19_18;
  assign nG_20_17 = nG_20_19 | (nP_20_19 & nG_18_17);
  assign nP_20_17 = nP_20_19 & nP_18_17;
  assign nG_19_16 = nG_19_18 | (nP_19_18 & nG_17_16);
  assign nP_19_16 = nP_19_18 & nP_17_16;
  assign nG_18_15 = nG_18_17 | (nP_18_17 & nG_16_15);
  assign nP_18_15 = nP_18_17 & nP_16_15;
  assign nG_17_14 = nG_17_16 | (nP_17_16 & nG_15_14);
  assign nP_17_14 = nP_17_16 & nP_15_14;
  assign nG_16_13 = nG_16_15 | (nP_16_15 & nG_14_13);
  assign nP_16_13 = nP_16_15 & nP_14_13;
  assign nG_15_12 = nG_15_14 | (nP_15_14 & nG_13_12);
  assign nP_15_12 = nP_15_14 & nP_13_12;
  assign nG_14_11 = nG_14_13 | (nP_14_13 & nG_12_11);
  assign nP_14_11 = nP_14_13 & nP_12_11;
  assign nG_13_10 = nG_13_12 | (nP_13_12 & nG_11_10);
  assign nP_13_10 = nP_13_12 & nP_11_10;
  assign nG_12_9 = nG_12_11 | (nP_12_11 & nG_10_9);
  assign nP_12_9 = nP_12_11 & nP_10_9;
  assign nG_11_8 = nG_11_10 | (nP_11_10 & nG_9_8);
  assign nP_11_8 = nP_11_10 & nP_9_8;
  assign nG_10_7 = nG_10_9 | (nP_10_9 & nG_8_7);
  assign nP_10_7 = nP_10_9 & nP_8_7;
  assign nG_9_6 = nG_9_8 | (nP_9_8 & nG_7_6);
  assign nP_9_6 = nP_9_8 & nP_7_6;
  assign nG_8_5 = nG_8_7 | (nP_8_7 & nG_6_5);
  assign nP_8_5 = nP_8_7 & nP_6_5;
  assign nG_7_4 = nG_7_6 | (nP_7_6 & nG_5_4);
  assign nP_7_4 = nP_7_6 & nP_5_4;
  assign nG_6_3 = nG_6_5 | (nP_6_5 & nG_4_3);
  assign nP_6_3 = nP_6_5 & nP_4_3;
  assign nG_5_2 = nG_5_4 | (nP_5_4 & nG_3_2);
  assign nP_5_2 = nP_5_4 & nP_3_2;
  assign nG_4_1 = nG_4_3 | (nP_4_3 & nG_2_1);
  assign nP_4_1 = nP_4_3 & nP_2_1;
  assign nG_3_0 = nG_3_2 | (nP_3_2 & nG_1_0);
  assign nP_3_0 = nP_3_2 & nP_1_0;
  assign nG_2_0 = nG_2_1 | (nP_2_1 & nG_0_0);
  assign nP_2_0 = nP_2_1 & nP_0_0;

  assign nG_63_56 = nG_63_60 | (nP_63_60 & nG_59_56);
  assign nP_63_56 = nP_63_60 & nP_59_56;
  assign nG_62_55 = nG_62_59 | (nP_62_59 & nG_58_55);
  assign nP_62_55 = nP_62_59 & nP_58_55;
  assign nG_61_54 = nG_61_58 | (nP_61_58 & nG_57_54);
  assign nP_61_54 = nP_61_58 & nP_57_54;
  assign nG_60_53 = nG_60_57 | (nP_60_57 & nG_56_53);
  assign nP_60_53 = nP_60_57 & nP_56_53;
  assign nG_59_52 = nG_59_56 | (nP_59_56 & nG_55_52);
  assign nP_59_52 = nP_59_56 & nP_55_52;
  assign nG_58_51 = nG_58_55 | (nP_58_55 & nG_54_51);
  assign nP_58_51 = nP_58_55 & nP_54_51;
  assign nG_57_50 = nG_57_54 | (nP_57_54 & nG_53_50);
  assign nP_57_50 = nP_57_54 & nP_53_50;
  assign nG_56_49 = nG_56_53 | (nP_56_53 & nG_52_49);
  assign nP_56_49 = nP_56_53 & nP_52_49;
  assign nG_55_48 = nG_55_52 | (nP_55_52 & nG_51_48);
  assign nP_55_48 = nP_55_52 & nP_51_48;
  assign nG_54_47 = nG_54_51 | (nP_54_51 & nG_50_47);
  assign nP_54_47 = nP_54_51 & nP_50_47;
  assign nG_53_46 = nG_53_50 | (nP_53_50 & nG_49_46);
  assign nP_53_46 = nP_53_50 & nP_49_46;
  assign nG_52_45 = nG_52_49 | (nP_52_49 & nG_48_45);
  assign nP_52_45 = nP_52_49 & nP_48_45;
  assign nG_51_44 = nG_51_48 | (nP_51_48 & nG_47_44);
  assign nP_51_44 = nP_51_48 & nP_47_44;
  assign nG_50_43 = nG_50_47 | (nP_50_47 & nG_46_43);
  assign nP_50_43 = nP_50_47 & nP_46_43;
  assign nG_49_42 = nG_49_46 | (nP_49_46 & nG_45_42);
  assign nP_49_42 = nP_49_46 & nP_45_42;
  assign nG_48_41 = nG_48_45 | (nP_48_45 & nG_44_41);
  assign nP_48_41 = nP_48_45 & nP_44_41;
  assign nG_47_40 = nG_47_44 | (nP_47_44 & nG_43_40);
  assign nP_47_40 = nP_47_44 & nP_43_40;
  assign nG_46_39 = nG_46_43 | (nP_46_43 & nG_42_39);
  assign nP_46_39 = nP_46_43 & nP_42_39;
  assign nG_45_38 = nG_45_42 | (nP_45_42 & nG_41_38);
  assign nP_45_38 = nP_45_42 & nP_41_38;
  assign nG_44_37 = nG_44_41 | (nP_44_41 & nG_40_37);
  assign nP_44_37 = nP_44_41 & nP_40_37;
  assign nG_43_36 = nG_43_40 | (nP_43_40 & nG_39_36);
  assign nP_43_36 = nP_43_40 & nP_39_36;
  assign nG_42_35 = nG_42_39 | (nP_42_39 & nG_38_35);
  assign nP_42_35 = nP_42_39 & nP_38_35;
  assign nG_41_34 = nG_41_38 | (nP_41_38 & nG_37_34);
  assign nP_41_34 = nP_41_38 & nP_37_34;
  assign nG_40_33 = nG_40_37 | (nP_40_37 & nG_36_33);
  assign nP_40_33 = nP_40_37 & nP_36_33;
  assign nG_39_32 = nG_39_36 | (nP_39_36 & nG_35_32);
  assign nP_39_32 = nP_39_36 & nP_35_32;
  assign nG_38_31 = nG_38_35 | (nP_38_35 & nG_34_31);
  assign nP_38_31 = nP_38_35 & nP_34_31;
  assign nG_37_30 = nG_37_34 | (nP_37_34 & nG_33_30);
  assign nP_37_30 = nP_37_34 & nP_33_30;
  assign nG_36_29 = nG_36_33 | (nP_36_33 & nG_32_29);
  assign nP_36_29 = nP_36_33 & nP_32_29;
  assign nG_35_28 = nG_35_32 | (nP_35_32 & nG_31_28);
  assign nP_35_28 = nP_35_32 & nP_31_28;
  assign nG_34_27 = nG_34_31 | (nP_34_31 & nG_30_27);
  assign nP_34_27 = nP_34_31 & nP_30_27;
  assign nG_33_26 = nG_33_30 | (nP_33_30 & nG_29_26);
  assign nP_33_26 = nP_33_30 & nP_29_26;
  assign nG_32_25 = nG_32_29 | (nP_32_29 & nG_28_25);
  assign nP_32_25 = nP_32_29 & nP_28_25;
  assign nG_31_24 = nG_31_28 | (nP_31_28 & nG_27_24);
  assign nP_31_24 = nP_31_28 & nP_27_24;
  assign nG_30_23 = nG_30_27 | (nP_30_27 & nG_26_23);
  assign nP_30_23 = nP_30_27 & nP_26_23;
  assign nG_29_22 = nG_29_26 | (nP_29_26 & nG_25_22);
  assign nP_29_22 = nP_29_26 & nP_25_22;
  assign nG_28_21 = nG_28_25 | (nP_28_25 & nG_24_21);
  assign nP_28_21 = nP_28_25 & nP_24_21;
  assign nG_27_20 = nG_27_24 | (nP_27_24 & nG_23_20);
  assign nP_27_20 = nP_27_24 & nP_23_20;
  assign nG_26_19 = nG_26_23 | (nP_26_23 & nG_22_19);
  assign nP_26_19 = nP_26_23 & nP_22_19;
  assign nG_25_18 = nG_25_22 | (nP_25_22 & nG_21_18);
  assign nP_25_18 = nP_25_22 & nP_21_18;
  assign nG_24_17 = nG_24_21 | (nP_24_21 & nG_20_17);
  assign nP_24_17 = nP_24_21 & nP_20_17;
  assign nG_23_16 = nG_23_20 | (nP_23_20 & nG_19_16);
  assign nP_23_16 = nP_23_20 & nP_19_16;
  assign nG_22_15 = nG_22_19 | (nP_22_19 & nG_18_15);
  assign nP_22_15 = nP_22_19 & nP_18_15;
  assign nG_21_14 = nG_21_18 | (nP_21_18 & nG_17_14);
  assign nP_21_14 = nP_21_18 & nP_17_14;
  assign nG_20_13 = nG_20_17 | (nP_20_17 & nG_16_13);
  assign nP_20_13 = nP_20_17 & nP_16_13;
  assign nG_19_12 = nG_19_16 | (nP_19_16 & nG_15_12);
  assign nP_19_12 = nP_19_16 & nP_15_12;
  assign nG_18_11 = nG_18_15 | (nP_18_15 & nG_14_11);
  assign nP_18_11 = nP_18_15 & nP_14_11;
  assign nG_17_10 = nG_17_14 | (nP_17_14 & nG_13_10);
  assign nP_17_10 = nP_17_14 & nP_13_10;
  assign nG_16_9 = nG_16_13 | (nP_16_13 & nG_12_9);
  assign nP_16_9 = nP_16_13 & nP_12_9;
  assign nG_15_8 = nG_15_12 | (nP_15_12 & nG_11_8);
  assign nP_15_8 = nP_15_12 & nP_11_8;
  assign nG_14_7 = nG_14_11 | (nP_14_11 & nG_10_7);
  assign nP_14_7 = nP_14_11 & nP_10_7;
  assign nG_13_6 = nG_13_10 | (nP_13_10 & nG_9_6);
  assign nP_13_6 = nP_13_10 & nP_9_6;
  assign nG_12_5 = nG_12_9 | (nP_12_9 & nG_8_5);
  assign nP_12_5 = nP_12_9 & nP_8_5;
  assign nG_11_4 = nG_11_8 | (nP_11_8 & nG_7_4);
  assign nP_11_4 = nP_11_8 & nP_7_4;
  assign nG_10_3 = nG_10_7 | (nP_10_7 & nG_6_3);
  assign nP_10_3 = nP_10_7 & nP_6_3;
  assign nG_9_2 = nG_9_6 | (nP_9_6 & nG_5_2);
  assign nP_9_2 = nP_9_6 & nP_5_2;
  assign nG_8_1 = nG_8_5 | (nP_8_5 & nG_4_1);
  assign nP_8_1 = nP_8_5 & nP_4_1;
  assign nG_7_0 = nG_7_4 | (nP_7_4 & nG_3_0);
  assign nP_7_0 = nP_7_4 & nP_3_0;
  assign nG_6_0 = nG_6_3 | (nP_6_3 & nG_2_0);
  assign nP_6_0 = nP_6_3 & nP_2_0;
  assign nG_5_0 = nG_5_2 | (nP_5_2 & nG_1_0);
  assign nP_5_0 = nP_5_2 & nP_1_0;
  assign nG_4_0 = nG_4_1 | (nP_4_1 & nG_0_0);
  assign nP_4_0 = nP_4_1 & nP_0_0;

  assign nG_63_48 = nG_63_56 | (nP_63_56 & nG_55_48);
  assign nP_63_48 = nP_63_56 & nP_55_48;
  assign nG_62_47 = nG_62_55 | (nP_62_55 & nG_54_47);
  assign nP_62_47 = nP_62_55 & nP_54_47;
  assign nG_61_46 = nG_61_54 | (nP_61_54 & nG_53_46);
  assign nP_61_46 = nP_61_54 & nP_53_46;
  assign nG_60_45 = nG_60_53 | (nP_60_53 & nG_52_45);
  assign nP_60_45 = nP_60_53 & nP_52_45;
  assign nG_59_44 = nG_59_52 | (nP_59_52 & nG_51_44);
  assign nP_59_44 = nP_59_52 & nP_51_44;
  assign nG_58_43 = nG_58_51 | (nP_58_51 & nG_50_43);
  assign nP_58_43 = nP_58_51 & nP_50_43;
  assign nG_57_42 = nG_57_50 | (nP_57_50 & nG_49_42);
  assign nP_57_42 = nP_57_50 & nP_49_42;
  assign nG_56_41 = nG_56_49 | (nP_56_49 & nG_48_41);
  assign nP_56_41 = nP_56_49 & nP_48_41;
  assign nG_55_40 = nG_55_48 | (nP_55_48 & nG_47_40);
  assign nP_55_40 = nP_55_48 & nP_47_40;
  assign nG_54_39 = nG_54_47 | (nP_54_47 & nG_46_39);
  assign nP_54_39 = nP_54_47 & nP_46_39;
  assign nG_53_38 = nG_53_46 | (nP_53_46 & nG_45_38);
  assign nP_53_38 = nP_53_46 & nP_45_38;
  assign nG_52_37 = nG_52_45 | (nP_52_45 & nG_44_37);
  assign nP_52_37 = nP_52_45 & nP_44_37;
  assign nG_51_36 = nG_51_44 | (nP_51_44 & nG_43_36);
  assign nP_51_36 = nP_51_44 & nP_43_36;
  assign nG_50_35 = nG_50_43 | (nP_50_43 & nG_42_35);
  assign nP_50_35 = nP_50_43 & nP_42_35;
  assign nG_49_34 = nG_49_42 | (nP_49_42 & nG_41_34);
  assign nP_49_34 = nP_49_42 & nP_41_34;
  assign nG_48_33 = nG_48_41 | (nP_48_41 & nG_40_33);
  assign nP_48_33 = nP_48_41 & nP_40_33;
  assign nG_47_32 = nG_47_40 | (nP_47_40 & nG_39_32);
  assign nP_47_32 = nP_47_40 & nP_39_32;
  assign nG_46_31 = nG_46_39 | (nP_46_39 & nG_38_31);
  assign nP_46_31 = nP_46_39 & nP_38_31;
  assign nG_45_30 = nG_45_38 | (nP_45_38 & nG_37_30);
  assign nP_45_30 = nP_45_38 & nP_37_30;
  assign nG_44_29 = nG_44_37 | (nP_44_37 & nG_36_29);
  assign nP_44_29 = nP_44_37 & nP_36_29;
  assign nG_43_28 = nG_43_36 | (nP_43_36 & nG_35_28);
  assign nP_43_28 = nP_43_36 & nP_35_28;
  assign nG_42_27 = nG_42_35 | (nP_42_35 & nG_34_27);
  assign nP_42_27 = nP_42_35 & nP_34_27;
  assign nG_41_26 = nG_41_34 | (nP_41_34 & nG_33_26);
  assign nP_41_26 = nP_41_34 & nP_33_26;
  assign nG_40_25 = nG_40_33 | (nP_40_33 & nG_32_25);
  assign nP_40_25 = nP_40_33 & nP_32_25;
  assign nG_39_24 = nG_39_32 | (nP_39_32 & nG_31_24);
  assign nP_39_24 = nP_39_32 & nP_31_24;
  assign nG_38_23 = nG_38_31 | (nP_38_31 & nG_30_23);
  assign nP_38_23 = nP_38_31 & nP_30_23;
  assign nG_37_22 = nG_37_30 | (nP_37_30 & nG_29_22);
  assign nP_37_22 = nP_37_30 & nP_29_22;
  assign nG_36_21 = nG_36_29 | (nP_36_29 & nG_28_21);
  assign nP_36_21 = nP_36_29 & nP_28_21;
  assign nG_35_20 = nG_35_28 | (nP_35_28 & nG_27_20);
  assign nP_35_20 = nP_35_28 & nP_27_20;
  assign nG_34_19 = nG_34_27 | (nP_34_27 & nG_26_19);
  assign nP_34_19 = nP_34_27 & nP_26_19;
  assign nG_33_18 = nG_33_26 | (nP_33_26 & nG_25_18);
  assign nP_33_18 = nP_33_26 & nP_25_18;
  assign nG_32_17 = nG_32_25 | (nP_32_25 & nG_24_17);
  assign nP_32_17 = nP_32_25 & nP_24_17;
  assign nG_31_16 = nG_31_24 | (nP_31_24 & nG_23_16);
  assign nP_31_16 = nP_31_24 & nP_23_16;
  assign nG_30_15 = nG_30_23 | (nP_30_23 & nG_22_15);
  assign nP_30_15 = nP_30_23 & nP_22_15;
  assign nG_29_14 = nG_29_22 | (nP_29_22 & nG_21_14);
  assign nP_29_14 = nP_29_22 & nP_21_14;
  assign nG_28_13 = nG_28_21 | (nP_28_21 & nG_20_13);
  assign nP_28_13 = nP_28_21 & nP_20_13;
  assign nG_27_12 = nG_27_20 | (nP_27_20 & nG_19_12);
  assign nP_27_12 = nP_27_20 & nP_19_12;
  assign nG_26_11 = nG_26_19 | (nP_26_19 & nG_18_11);
  assign nP_26_11 = nP_26_19 & nP_18_11;
  assign nG_25_10 = nG_25_18 | (nP_25_18 & nG_17_10);
  assign nP_25_10 = nP_25_18 & nP_17_10;
  assign nG_24_9 = nG_24_17 | (nP_24_17 & nG_16_9);
  assign nP_24_9 = nP_24_17 & nP_16_9;
  assign nG_23_8 = nG_23_16 | (nP_23_16 & nG_15_8);
  assign nP_23_8 = nP_23_16 & nP_15_8;
  assign nG_22_7 = nG_22_15 | (nP_22_15 & nG_14_7);
  assign nP_22_7 = nP_22_15 & nP_14_7;
  assign nG_21_6 = nG_21_14 | (nP_21_14 & nG_13_6);
  assign nP_21_6 = nP_21_14 & nP_13_6;
  assign nG_20_5 = nG_20_13 | (nP_20_13 & nG_12_5);
  assign nP_20_5 = nP_20_13 & nP_12_5;
  assign nG_19_4 = nG_19_12 | (nP_19_12 & nG_11_4);
  assign nP_19_4 = nP_19_12 & nP_11_4;
  assign nG_18_3 = nG_18_11 | (nP_18_11 & nG_10_3);
  assign nP_18_3 = nP_18_11 & nP_10_3;
  assign nG_17_2 = nG_17_10 | (nP_17_10 & nG_9_2);
  assign nP_17_2 = nP_17_10 & nP_9_2;
  assign nG_16_1 = nG_16_9 | (nP_16_9 & nG_8_1);
  assign nP_16_1 = nP_16_9 & nP_8_1;
  assign nG_15_0 = nG_15_8 | (nP_15_8 & nG_7_0);
  assign nP_15_0 = nP_15_8 & nP_7_0;
  assign nG_14_0 = nG_14_7 | (nP_14_7 & nG_6_0);
  assign nP_14_0 = nP_14_7 & nP_6_0;
  assign nG_13_0 = nG_13_6 | (nP_13_6 & nG_5_0);
  assign nP_13_0 = nP_13_6 & nP_5_0;
  assign nG_12_0 = nG_12_5 | (nP_12_5 & nG_4_0);
  assign nP_12_0 = nP_12_5 & nP_4_0;
  assign nG_11_0 = nG_11_4 | (nP_11_4 & nG_3_0);
  assign nP_11_0 = nP_11_4 & nP_3_0;
  assign nG_10_0 = nG_10_3 | (nP_10_3 & nG_2_0);
  assign nP_10_0 = nP_10_3 & nP_2_0;
  assign nG_9_0 = nG_9_2 | (nP_9_2 & nG_1_0);
  assign nP_9_0 = nP_9_2 & nP_1_0;
  assign nG_8_0 = nG_8_1 | (nP_8_1 & nG_0_0);
  assign nP_8_0 = nP_8_1 & nP_0_0;

  assign nG_63_32 = nG_63_48 | (nP_63_48 & nG_47_32);
  assign nP_63_32 = nP_63_48 & nP_47_32;
  assign nG_62_31 = nG_62_47 | (nP_62_47 & nG_46_31);
  assign nP_62_31 = nP_62_47 & nP_46_31;
  assign nG_61_30 = nG_61_46 | (nP_61_46 & nG_45_30);
  assign nP_61_30 = nP_61_46 & nP_45_30;
  assign nG_60_29 = nG_60_45 | (nP_60_45 & nG_44_29);
  assign nP_60_29 = nP_60_45 & nP_44_29;
  assign nG_59_28 = nG_59_44 | (nP_59_44 & nG_43_28);
  assign nP_59_28 = nP_59_44 & nP_43_28;
  assign nG_58_27 = nG_58_43 | (nP_58_43 & nG_42_27);
  assign nP_58_27 = nP_58_43 & nP_42_27;
  assign nG_57_26 = nG_57_42 | (nP_57_42 & nG_41_26);
  assign nP_57_26 = nP_57_42 & nP_41_26;
  assign nG_56_25 = nG_56_41 | (nP_56_41 & nG_40_25);
  assign nP_56_25 = nP_56_41 & nP_40_25;
  assign nG_55_24 = nG_55_40 | (nP_55_40 & nG_39_24);
  assign nP_55_24 = nP_55_40 & nP_39_24;
  assign nG_54_23 = nG_54_39 | (nP_54_39 & nG_38_23);
  assign nP_54_23 = nP_54_39 & nP_38_23;
  assign nG_53_22 = nG_53_38 | (nP_53_38 & nG_37_22);
  assign nP_53_22 = nP_53_38 & nP_37_22;
  assign nG_52_21 = nG_52_37 | (nP_52_37 & nG_36_21);
  assign nP_52_21 = nP_52_37 & nP_36_21;
  assign nG_51_20 = nG_51_36 | (nP_51_36 & nG_35_20);
  assign nP_51_20 = nP_51_36 & nP_35_20;
  assign nG_50_19 = nG_50_35 | (nP_50_35 & nG_34_19);
  assign nP_50_19 = nP_50_35 & nP_34_19;
  assign nG_49_18 = nG_49_34 | (nP_49_34 & nG_33_18);
  assign nP_49_18 = nP_49_34 & nP_33_18;
  assign nG_48_17 = nG_48_33 | (nP_48_33 & nG_32_17);
  assign nP_48_17 = nP_48_33 & nP_32_17;
  assign nG_47_16 = nG_47_32 | (nP_47_32 & nG_31_16);
  assign nP_47_16 = nP_47_32 & nP_31_16;
  assign nG_46_15 = nG_46_31 | (nP_46_31 & nG_30_15);
  assign nP_46_15 = nP_46_31 & nP_30_15;
  assign nG_45_14 = nG_45_30 | (nP_45_30 & nG_29_14);
  assign nP_45_14 = nP_45_30 & nP_29_14;
  assign nG_44_13 = nG_44_29 | (nP_44_29 & nG_28_13);
  assign nP_44_13 = nP_44_29 & nP_28_13;
  assign nG_43_12 = nG_43_28 | (nP_43_28 & nG_27_12);
  assign nP_43_12 = nP_43_28 & nP_27_12;
  assign nG_42_11 = nG_42_27 | (nP_42_27 & nG_26_11);
  assign nP_42_11 = nP_42_27 & nP_26_11;
  assign nG_41_10 = nG_41_26 | (nP_41_26 & nG_25_10);
  assign nP_41_10 = nP_41_26 & nP_25_10;
  assign nG_40_9 = nG_40_25 | (nP_40_25 & nG_24_9);
  assign nP_40_9 = nP_40_25 & nP_24_9;
  assign nG_39_8 = nG_39_24 | (nP_39_24 & nG_23_8);
  assign nP_39_8 = nP_39_24 & nP_23_8;
  assign nG_38_7 = nG_38_23 | (nP_38_23 & nG_22_7);
  assign nP_38_7 = nP_38_23 & nP_22_7;
  assign nG_37_6 = nG_37_22 | (nP_37_22 & nG_21_6);
  assign nP_37_6 = nP_37_22 & nP_21_6;
  assign nG_36_5 = nG_36_21 | (nP_36_21 & nG_20_5);
  assign nP_36_5 = nP_36_21 & nP_20_5;
  assign nG_35_4 = nG_35_20 | (nP_35_20 & nG_19_4);
  assign nP_35_4 = nP_35_20 & nP_19_4;
  assign nG_34_3 = nG_34_19 | (nP_34_19 & nG_18_3);
  assign nP_34_3 = nP_34_19 & nP_18_3;
  assign nG_33_2 = nG_33_18 | (nP_33_18 & nG_17_2);
  assign nP_33_2 = nP_33_18 & nP_17_2;
  assign nG_32_1 = nG_32_17 | (nP_32_17 & nG_16_1);
  assign nP_32_1 = nP_32_17 & nP_16_1;
  assign nG_31_0 = nG_31_16 | (nP_31_16 & nG_15_0);
  assign nP_31_0 = nP_31_16 & nP_15_0;
  assign nG_30_0 = nG_30_15 | (nP_30_15 & nG_14_0);
  assign nP_30_0 = nP_30_15 & nP_14_0;
  assign nG_29_0 = nG_29_14 | (nP_29_14 & nG_13_0);
  assign nP_29_0 = nP_29_14 & nP_13_0;
  assign nG_28_0 = nG_28_13 | (nP_28_13 & nG_12_0);
  assign nP_28_0 = nP_28_13 & nP_12_0;
  assign nG_27_0 = nG_27_12 | (nP_27_12 & nG_11_0);
  assign nP_27_0 = nP_27_12 & nP_11_0;
  assign nG_26_0 = nG_26_11 | (nP_26_11 & nG_10_0);
  assign nP_26_0 = nP_26_11 & nP_10_0;
  assign nG_25_0 = nG_25_10 | (nP_25_10 & nG_9_0);
  assign nP_25_0 = nP_25_10 & nP_9_0;
  assign nG_24_0 = nG_24_9 | (nP_24_9 & nG_8_0);
  assign nP_24_0 = nP_24_9 & nP_8_0;
  assign nG_23_0 = nG_23_8 | (nP_23_8 & nG_7_0);
  assign nP_23_0 = nP_23_8 & nP_7_0;
  assign nG_22_0 = nG_22_7 | (nP_22_7 & nG_6_0);
  assign nP_22_0 = nP_22_7 & nP_6_0;
  assign nG_21_0 = nG_21_6 | (nP_21_6 & nG_5_0);
  assign nP_21_0 = nP_21_6 & nP_5_0;
  assign nG_20_0 = nG_20_5 | (nP_20_5 & nG_4_0);
  assign nP_20_0 = nP_20_5 & nP_4_0;
  assign nG_19_0 = nG_19_4 | (nP_19_4 & nG_3_0);
  assign nP_19_0 = nP_19_4 & nP_3_0;
  assign nG_18_0 = nG_18_3 | (nP_18_3 & nG_2_0);
  assign nP_18_0 = nP_18_3 & nP_2_0;
  assign nG_17_0 = nG_17_2 | (nP_17_2 & nG_1_0);
  assign nP_17_0 = nP_17_2 & nP_1_0;
  assign nG_16_0 = nG_16_1 | (nP_16_1 & nG_0_0);
  assign nP_16_0 = nP_16_1 & nP_0_0;

  assign nG_63_0 = nG_63_32 | (nP_63_32 & nG_31_0);
  assign nP_63_0 = nP_63_32 & nP_31_0;
  assign nG_62_0 = nG_62_31 | (nP_62_31 & nG_30_0);
  assign nP_62_0 = nP_62_31 & nP_30_0;
  assign nG_61_0 = nG_61_30 | (nP_61_30 & nG_29_0);
  assign nP_61_0 = nP_61_30 & nP_29_0;
  assign nG_60_0 = nG_60_29 | (nP_60_29 & nG_28_0);
  assign nP_60_0 = nP_60_29 & nP_28_0;
  assign nG_59_0 = nG_59_28 | (nP_59_28 & nG_27_0);
  assign nP_59_0 = nP_59_28 & nP_27_0;
  assign nG_58_0 = nG_58_27 | (nP_58_27 & nG_26_0);
  assign nP_58_0 = nP_58_27 & nP_26_0;
  assign nG_57_0 = nG_57_26 | (nP_57_26 & nG_25_0);
  assign nP_57_0 = nP_57_26 & nP_25_0;
  assign nG_56_0 = nG_56_25 | (nP_56_25 & nG_24_0);
  assign nP_56_0 = nP_56_25 & nP_24_0;
  assign nG_55_0 = nG_55_24 | (nP_55_24 & nG_23_0);
  assign nP_55_0 = nP_55_24 & nP_23_0;
  assign nG_54_0 = nG_54_23 | (nP_54_23 & nG_22_0);
  assign nP_54_0 = nP_54_23 & nP_22_0;
  assign nG_53_0 = nG_53_22 | (nP_53_22 & nG_21_0);
  assign nP_53_0 = nP_53_22 & nP_21_0;
  assign nG_52_0 = nG_52_21 | (nP_52_21 & nG_20_0);
  assign nP_52_0 = nP_52_21 & nP_20_0;
  assign nG_51_0 = nG_51_20 | (nP_51_20 & nG_19_0);
  assign nP_51_0 = nP_51_20 & nP_19_0;
  assign nG_50_0 = nG_50_19 | (nP_50_19 & nG_18_0);
  assign nP_50_0 = nP_50_19 & nP_18_0;
  assign nG_49_0 = nG_49_18 | (nP_49_18 & nG_17_0);
  assign nP_49_0 = nP_49_18 & nP_17_0;
  assign nG_48_0 = nG_48_17 | (nP_48_17 & nG_16_0);
  assign nP_48_0 = nP_48_17 & nP_16_0;
  assign nG_47_0 = nG_47_16 | (nP_47_16 & nG_15_0);
  assign nP_47_0 = nP_47_16 & nP_15_0;
  assign nG_46_0 = nG_46_15 | (nP_46_15 & nG_14_0);
  assign nP_46_0 = nP_46_15 & nP_14_0;
  assign nG_45_0 = nG_45_14 | (nP_45_14 & nG_13_0);
  assign nP_45_0 = nP_45_14 & nP_13_0;
  assign nG_44_0 = nG_44_13 | (nP_44_13 & nG_12_0);
  assign nP_44_0 = nP_44_13 & nP_12_0;
  assign nG_43_0 = nG_43_12 | (nP_43_12 & nG_11_0);
  assign nP_43_0 = nP_43_12 & nP_11_0;
  assign nG_42_0 = nG_42_11 | (nP_42_11 & nG_10_0);
  assign nP_42_0 = nP_42_11 & nP_10_0;
  assign nG_41_0 = nG_41_10 | (nP_41_10 & nG_9_0);
  assign nP_41_0 = nP_41_10 & nP_9_0;
  assign nG_40_0 = nG_40_9 | (nP_40_9 & nG_8_0);
  assign nP_40_0 = nP_40_9 & nP_8_0;
  assign nG_39_0 = nG_39_8 | (nP_39_8 & nG_7_0);
  assign nP_39_0 = nP_39_8 & nP_7_0;
  assign nG_38_0 = nG_38_7 | (nP_38_7 & nG_6_0);
  assign nP_38_0 = nP_38_7 & nP_6_0;
  assign nG_37_0 = nG_37_6 | (nP_37_6 & nG_5_0);
  assign nP_37_0 = nP_37_6 & nP_5_0;
  assign nG_36_0 = nG_36_5 | (nP_36_5 & nG_4_0);
  assign nP_36_0 = nP_36_5 & nP_4_0;
  assign nG_35_0 = nG_35_4 | (nP_35_4 & nG_3_0);
  assign nP_35_0 = nP_35_4 & nP_3_0;
  assign nG_34_0 = nG_34_3 | (nP_34_3 & nG_2_0);
  assign nP_34_0 = nP_34_3 & nP_2_0;
  assign nG_33_0 = nG_33_2 | (nP_33_2 & nG_1_0);
  assign nP_33_0 = nP_33_2 & nP_1_0;
  assign nG_32_0 = nG_32_1 | (nP_32_1 & nG_0_0);
  assign nP_32_0 = nP_32_1 & nP_0_0;

  assign nC_0 = in_CI;
  assign nC_1 = nG_0_0 | (nP_0_0 & in_CI);
  assign nC_2 = nG_1_0 | (nP_1_0 & in_CI);
  assign nC_3 = nG_2_0 | (nP_2_0 & in_CI);
  assign nC_4 = nG_3_0 | (nP_3_0 & in_CI);
  assign nC_5 = nG_4_0 | (nP_4_0 & in_CI);
  assign nC_6 = nG_5_0 | (nP_5_0 & in_CI);
  assign nC_7 = nG_6_0 | (nP_6_0 & in_CI);
  assign nC_8 = nG_7_0 | (nP_7_0 & in_CI);
  assign nC_9 = nG_8_0 | (nP_8_0 & in_CI);
  assign nC_10 = nG_9_0 | (nP_9_0 & in_CI);
  assign nC_11 = nG_10_0 | (nP_10_0 & in_CI);
  assign nC_12 = nG_11_0 | (nP_11_0 & in_CI);
  assign nC_13 = nG_12_0 | (nP_12_0 & in_CI);
  assign nC_14 = nG_13_0 | (nP_13_0 & in_CI);
  assign nC_15 = nG_14_0 | (nP_14_0 & in_CI);
  assign nC_16 = nG_15_0 | (nP_15_0 & in_CI);
  assign nC_17 = nG_16_0 | (nP_16_0 & in_CI);
  assign nC_18 = nG_17_0 | (nP_17_0 & in_CI);
  assign nC_19 = nG_18_0 | (nP_18_0 & in_CI);
  assign nC_20 = nG_19_0 | (nP_19_0 & in_CI);
  assign nC_21 = nG_20_0 | (nP_20_0 & in_CI);
  assign nC_22 = nG_21_0 | (nP_21_0 & in_CI);
  assign nC_23 = nG_22_0 | (nP_22_0 & in_CI);
  assign nC_24 = nG_23_0 | (nP_23_0 & in_CI);
  assign nC_25 = nG_24_0 | (nP_24_0 & in_CI);
  assign nC_26 = nG_25_0 | (nP_25_0 & in_CI);
  assign nC_27 = nG_26_0 | (nP_26_0 & in_CI);
  assign nC_28 = nG_27_0 | (nP_27_0 & in_CI);
  assign nC_29 = nG_28_0 | (nP_28_0 & in_CI);
  assign nC_30 = nG_29_0 | (nP_29_0 & in_CI);
  assign nC_31 = nG_30_0 | (nP_30_0 & in_CI);
  assign nC_32 = nG_31_0 | (nP_31_0 & in_CI);
  assign nC_33 = nG_32_0 | (nP_32_0 & in_CI);
  assign nC_34 = nG_33_0 | (nP_33_0 & in_CI);
  assign nC_35 = nG_34_0 | (nP_34_0 & in_CI);
  assign nC_36 = nG_35_0 | (nP_35_0 & in_CI);
  assign nC_37 = nG_36_0 | (nP_36_0 & in_CI);
  assign nC_38 = nG_37_0 | (nP_37_0 & in_CI);
  assign nC_39 = nG_38_0 | (nP_38_0 & in_CI);
  assign nC_40 = nG_39_0 | (nP_39_0 & in_CI);
  assign nC_41 = nG_40_0 | (nP_40_0 & in_CI);
  assign nC_42 = nG_41_0 | (nP_41_0 & in_CI);
  assign nC_43 = nG_42_0 | (nP_42_0 & in_CI);
  assign nC_44 = nG_43_0 | (nP_43_0 & in_CI);
  assign nC_45 = nG_44_0 | (nP_44_0 & in_CI);
  assign nC_46 = nG_45_0 | (nP_45_0 & in_CI);
  assign nC_47 = nG_46_0 | (nP_46_0 & in_CI);
  assign nC_48 = nG_47_0 | (nP_47_0 & in_CI);
  assign nC_49 = nG_48_0 | (nP_48_0 & in_CI);
  assign nC_50 = nG_49_0 | (nP_49_0 & in_CI);
  assign nC_51 = nG_50_0 | (nP_50_0 & in_CI);
  assign nC_52 = nG_51_0 | (nP_51_0 & in_CI);
  assign nC_53 = nG_52_0 | (nP_52_0 & in_CI);
  assign nC_54 = nG_53_0 | (nP_53_0 & in_CI);
  assign nC_55 = nG_54_0 | (nP_54_0 & in_CI);
  assign nC_56 = nG_55_0 | (nP_55_0 & in_CI);
  assign nC_57 = nG_56_0 | (nP_56_0 & in_CI);
  assign nC_58 = nG_57_0 | (nP_57_0 & in_CI);
  assign nC_59 = nG_58_0 | (nP_58_0 & in_CI);
  assign nC_60 = nG_59_0 | (nP_59_0 & in_CI);
  assign nC_61 = nG_60_0 | (nP_60_0 & in_CI);
  assign nC_62 = nG_61_0 | (nP_61_0 & in_CI);
  assign nC_63 = nG_62_0 | (nP_62_0 & in_CI);

  assign out_S[0] = nP_0_0 ^ nC_0;
  assign out_S[1] = nP_1_1 ^ nC_1;
  assign out_S[2] = nP_2_2 ^ nC_2;
  assign out_S[3] = nP_3_3 ^ nC_3;
  assign out_S[4] = nP_4_4 ^ nC_4;
  assign out_S[5] = nP_5_5 ^ nC_5;
  assign out_S[6] = nP_6_6 ^ nC_6;
  assign out_S[7] = nP_7_7 ^ nC_7;
  assign out_S[8] = nP_8_8 ^ nC_8;
  assign out_S[9] = nP_9_9 ^ nC_9;
  assign out_S[10] = nP_10_10 ^ nC_10;
  assign out_S[11] = nP_11_11 ^ nC_11;
  assign out_S[12] = nP_12_12 ^ nC_12;
  assign out_S[13] = nP_13_13 ^ nC_13;
  assign out_S[14] = nP_14_14 ^ nC_14;
  assign out_S[15] = nP_15_15 ^ nC_15;
  assign out_S[16] = nP_16_16 ^ nC_16;
  assign out_S[17] = nP_17_17 ^ nC_17;
  assign out_S[18] = nP_18_18 ^ nC_18;
  assign out_S[19] = nP_19_19 ^ nC_19;
  assign out_S[20] = nP_20_20 ^ nC_20;
  assign out_S[21] = nP_21_21 ^ nC_21;
  assign out_S[22] = nP_22_22 ^ nC_22;
  assign out_S[23] = nP_23_23 ^ nC_23;
  assign out_S[24] = nP_24_24 ^ nC_24;
  assign out_S[25] = nP_25_25 ^ nC_25;
  assign out_S[26] = nP_26_26 ^ nC_26;
  assign out_S[27] = nP_27_27 ^ nC_27;
  assign out_S[28] = nP_28_28 ^ nC_28;
  assign out_S[29] = nP_29_29 ^ nC_29;
  assign out_S[30] = nP_30_30 ^ nC_30;
  assign out_S[31] = nP_31_31 ^ nC_31;
  assign out_S[32] = nP_32_32 ^ nC_32;
  assign out_S[33] = nP_33_33 ^ nC_33;
  assign out_S[34] = nP_34_34 ^ nC_34;
  assign out_S[35] = nP_35_35 ^ nC_35;
  assign out_S[36] = nP_36_36 ^ nC_36;
  assign out_S[37] = nP_37_37 ^ nC_37;
  assign out_S[38] = nP_38_38 ^ nC_38;
  assign out_S[39] = nP_39_39 ^ nC_39;
  assign out_S[40] = nP_40_40 ^ nC_40;
  assign out_S[41] = nP_41_41 ^ nC_41;
  assign out_S[42] = nP_42_42 ^ nC_42;
  assign out_S[43] = nP_43_43 ^ nC_43;
  assign out_S[44] = nP_44_44 ^ nC_44;
  assign out_S[45] = nP_45_45 ^ nC_45;
  assign out_S[46] = nP_46_46 ^ nC_46;
  assign out_S[47] = nP_47_47 ^ nC_47;
  assign out_S[48] = nP_48_48 ^ nC_48;
  assign out_S[49] = nP_49_49 ^ nC_49;
  assign out_S[50] = nP_50_50 ^ nC_50;
  assign out_S[51] = nP_51_51 ^ nC_51;
  assign out_S[52] = nP_52_52 ^ nC_52;
  assign out_S[53] = nP_53_53 ^ nC_53;
  assign out_S[54] = nP_54_54 ^ nC_54;
  assign out_S[55] = nP_55_55 ^ nC_55;
  assign out_S[56] = nP_56_56 ^ nC_56;
  assign out_S[57] = nP_57_57 ^ nC_57;
  assign out_S[58] = nP_58_58 ^ nC_58;
  assign out_S[59] = nP_59_59 ^ nC_59;
  assign out_S[60] = nP_60_60 ^ nC_60;
  assign out_S[61] = nP_61_61 ^ nC_61;
  assign out_S[62] = nP_62_62 ^ nC_62;
  assign out_S[63] = nP_63_63 ^ nC_63;
  assign out_CO = nG_63_0 | (nP_63_0 & in_CI);
endmodule

