/net/ugrads/jtschir1/pvt/ee434/lab3/lib/lef/NangateOpenCellLibrary.lef