module VFA (in_A, in_B, in_CI, out_S, out_CO);
  input in_A, in_B, in_CI;
  output out_S, out_CO;

  assign out_S = in_A ^ in_B ^ in_CI;
  assign out_CO = (in_A & in_B) | (in_B & in_CI) | (in_CI & in_A);
endmodule



module VRCA_256 (in_A, in_B, in_CI, out_S, out_CO);
  input [255:0] in_A, in_B;
  input in_CI;
  output [255:0] out_S;
  output out_CO;

  VFA U0 (.in_A(in_A[0]), .in_B(in_B[0]), .in_CI(in_CI), .out_S(out_S[0]), .out_CO(nC1));
  VFA U1 (.in_A(in_A[1]), .in_B(in_B[1]), .in_CI(nC1), .out_S(out_S[1]), .out_CO(nC2));
  VFA U2 (.in_A(in_A[2]), .in_B(in_B[2]), .in_CI(nC2), .out_S(out_S[2]), .out_CO(nC3));
  VFA U3 (.in_A(in_A[3]), .in_B(in_B[3]), .in_CI(nC3), .out_S(out_S[3]), .out_CO(nC4));
  VFA U4 (.in_A(in_A[4]), .in_B(in_B[4]), .in_CI(nC4), .out_S(out_S[4]), .out_CO(nC5));
  VFA U5 (.in_A(in_A[5]), .in_B(in_B[5]), .in_CI(nC5), .out_S(out_S[5]), .out_CO(nC6));
  VFA U6 (.in_A(in_A[6]), .in_B(in_B[6]), .in_CI(nC6), .out_S(out_S[6]), .out_CO(nC7));
  VFA U7 (.in_A(in_A[7]), .in_B(in_B[7]), .in_CI(nC7), .out_S(out_S[7]), .out_CO(nC8));
  VFA U8 (.in_A(in_A[8]), .in_B(in_B[8]), .in_CI(nC8), .out_S(out_S[8]), .out_CO(nC9));
  VFA U9 (.in_A(in_A[9]), .in_B(in_B[9]), .in_CI(nC9), .out_S(out_S[9]), .out_CO(nC10));
  VFA U10 (.in_A(in_A[10]), .in_B(in_B[10]), .in_CI(nC10), .out_S(out_S[10]), .out_CO(nC11));
  VFA U11 (.in_A(in_A[11]), .in_B(in_B[11]), .in_CI(nC11), .out_S(out_S[11]), .out_CO(nC12));
  VFA U12 (.in_A(in_A[12]), .in_B(in_B[12]), .in_CI(nC12), .out_S(out_S[12]), .out_CO(nC13));
  VFA U13 (.in_A(in_A[13]), .in_B(in_B[13]), .in_CI(nC13), .out_S(out_S[13]), .out_CO(nC14));
  VFA U14 (.in_A(in_A[14]), .in_B(in_B[14]), .in_CI(nC14), .out_S(out_S[14]), .out_CO(nC15));
  VFA U15 (.in_A(in_A[15]), .in_B(in_B[15]), .in_CI(nC15), .out_S(out_S[15]), .out_CO(nC16));
  VFA U16 (.in_A(in_A[16]), .in_B(in_B[16]), .in_CI(nC16), .out_S(out_S[16]), .out_CO(nC17));
  VFA U17 (.in_A(in_A[17]), .in_B(in_B[17]), .in_CI(nC17), .out_S(out_S[17]), .out_CO(nC18));
  VFA U18 (.in_A(in_A[18]), .in_B(in_B[18]), .in_CI(nC18), .out_S(out_S[18]), .out_CO(nC19));
  VFA U19 (.in_A(in_A[19]), .in_B(in_B[19]), .in_CI(nC19), .out_S(out_S[19]), .out_CO(nC20));
  VFA U20 (.in_A(in_A[20]), .in_B(in_B[20]), .in_CI(nC20), .out_S(out_S[20]), .out_CO(nC21));
  VFA U21 (.in_A(in_A[21]), .in_B(in_B[21]), .in_CI(nC21), .out_S(out_S[21]), .out_CO(nC22));
  VFA U22 (.in_A(in_A[22]), .in_B(in_B[22]), .in_CI(nC22), .out_S(out_S[22]), .out_CO(nC23));
  VFA U23 (.in_A(in_A[23]), .in_B(in_B[23]), .in_CI(nC23), .out_S(out_S[23]), .out_CO(nC24));
  VFA U24 (.in_A(in_A[24]), .in_B(in_B[24]), .in_CI(nC24), .out_S(out_S[24]), .out_CO(nC25));
  VFA U25 (.in_A(in_A[25]), .in_B(in_B[25]), .in_CI(nC25), .out_S(out_S[25]), .out_CO(nC26));
  VFA U26 (.in_A(in_A[26]), .in_B(in_B[26]), .in_CI(nC26), .out_S(out_S[26]), .out_CO(nC27));
  VFA U27 (.in_A(in_A[27]), .in_B(in_B[27]), .in_CI(nC27), .out_S(out_S[27]), .out_CO(nC28));
  VFA U28 (.in_A(in_A[28]), .in_B(in_B[28]), .in_CI(nC28), .out_S(out_S[28]), .out_CO(nC29));
  VFA U29 (.in_A(in_A[29]), .in_B(in_B[29]), .in_CI(nC29), .out_S(out_S[29]), .out_CO(nC30));
  VFA U30 (.in_A(in_A[30]), .in_B(in_B[30]), .in_CI(nC30), .out_S(out_S[30]), .out_CO(nC31));
  VFA U31 (.in_A(in_A[31]), .in_B(in_B[31]), .in_CI(nC31), .out_S(out_S[31]), .out_CO(nC32));
  VFA U32 (.in_A(in_A[32]), .in_B(in_B[32]), .in_CI(nC32), .out_S(out_S[32]), .out_CO(nC33));
  VFA U33 (.in_A(in_A[33]), .in_B(in_B[33]), .in_CI(nC33), .out_S(out_S[33]), .out_CO(nC34));
  VFA U34 (.in_A(in_A[34]), .in_B(in_B[34]), .in_CI(nC34), .out_S(out_S[34]), .out_CO(nC35));
  VFA U35 (.in_A(in_A[35]), .in_B(in_B[35]), .in_CI(nC35), .out_S(out_S[35]), .out_CO(nC36));
  VFA U36 (.in_A(in_A[36]), .in_B(in_B[36]), .in_CI(nC36), .out_S(out_S[36]), .out_CO(nC37));
  VFA U37 (.in_A(in_A[37]), .in_B(in_B[37]), .in_CI(nC37), .out_S(out_S[37]), .out_CO(nC38));
  VFA U38 (.in_A(in_A[38]), .in_B(in_B[38]), .in_CI(nC38), .out_S(out_S[38]), .out_CO(nC39));
  VFA U39 (.in_A(in_A[39]), .in_B(in_B[39]), .in_CI(nC39), .out_S(out_S[39]), .out_CO(nC40));
  VFA U40 (.in_A(in_A[40]), .in_B(in_B[40]), .in_CI(nC40), .out_S(out_S[40]), .out_CO(nC41));
  VFA U41 (.in_A(in_A[41]), .in_B(in_B[41]), .in_CI(nC41), .out_S(out_S[41]), .out_CO(nC42));
  VFA U42 (.in_A(in_A[42]), .in_B(in_B[42]), .in_CI(nC42), .out_S(out_S[42]), .out_CO(nC43));
  VFA U43 (.in_A(in_A[43]), .in_B(in_B[43]), .in_CI(nC43), .out_S(out_S[43]), .out_CO(nC44));
  VFA U44 (.in_A(in_A[44]), .in_B(in_B[44]), .in_CI(nC44), .out_S(out_S[44]), .out_CO(nC45));
  VFA U45 (.in_A(in_A[45]), .in_B(in_B[45]), .in_CI(nC45), .out_S(out_S[45]), .out_CO(nC46));
  VFA U46 (.in_A(in_A[46]), .in_B(in_B[46]), .in_CI(nC46), .out_S(out_S[46]), .out_CO(nC47));
  VFA U47 (.in_A(in_A[47]), .in_B(in_B[47]), .in_CI(nC47), .out_S(out_S[47]), .out_CO(nC48));
  VFA U48 (.in_A(in_A[48]), .in_B(in_B[48]), .in_CI(nC48), .out_S(out_S[48]), .out_CO(nC49));
  VFA U49 (.in_A(in_A[49]), .in_B(in_B[49]), .in_CI(nC49), .out_S(out_S[49]), .out_CO(nC50));
  VFA U50 (.in_A(in_A[50]), .in_B(in_B[50]), .in_CI(nC50), .out_S(out_S[50]), .out_CO(nC51));
  VFA U51 (.in_A(in_A[51]), .in_B(in_B[51]), .in_CI(nC51), .out_S(out_S[51]), .out_CO(nC52));
  VFA U52 (.in_A(in_A[52]), .in_B(in_B[52]), .in_CI(nC52), .out_S(out_S[52]), .out_CO(nC53));
  VFA U53 (.in_A(in_A[53]), .in_B(in_B[53]), .in_CI(nC53), .out_S(out_S[53]), .out_CO(nC54));
  VFA U54 (.in_A(in_A[54]), .in_B(in_B[54]), .in_CI(nC54), .out_S(out_S[54]), .out_CO(nC55));
  VFA U55 (.in_A(in_A[55]), .in_B(in_B[55]), .in_CI(nC55), .out_S(out_S[55]), .out_CO(nC56));
  VFA U56 (.in_A(in_A[56]), .in_B(in_B[56]), .in_CI(nC56), .out_S(out_S[56]), .out_CO(nC57));
  VFA U57 (.in_A(in_A[57]), .in_B(in_B[57]), .in_CI(nC57), .out_S(out_S[57]), .out_CO(nC58));
  VFA U58 (.in_A(in_A[58]), .in_B(in_B[58]), .in_CI(nC58), .out_S(out_S[58]), .out_CO(nC59));
  VFA U59 (.in_A(in_A[59]), .in_B(in_B[59]), .in_CI(nC59), .out_S(out_S[59]), .out_CO(nC60));
  VFA U60 (.in_A(in_A[60]), .in_B(in_B[60]), .in_CI(nC60), .out_S(out_S[60]), .out_CO(nC61));
  VFA U61 (.in_A(in_A[61]), .in_B(in_B[61]), .in_CI(nC61), .out_S(out_S[61]), .out_CO(nC62));
  VFA U62 (.in_A(in_A[62]), .in_B(in_B[62]), .in_CI(nC62), .out_S(out_S[62]), .out_CO(nC63));
  VFA U63 (.in_A(in_A[63]), .in_B(in_B[63]), .in_CI(nC63), .out_S(out_S[63]), .out_CO(nC64));
  VFA U64 (.in_A(in_A[64]), .in_B(in_B[64]), .in_CI(nC64), .out_S(out_S[64]), .out_CO(nC65));
  VFA U65 (.in_A(in_A[65]), .in_B(in_B[65]), .in_CI(nC65), .out_S(out_S[65]), .out_CO(nC66));
  VFA U66 (.in_A(in_A[66]), .in_B(in_B[66]), .in_CI(nC66), .out_S(out_S[66]), .out_CO(nC67));
  VFA U67 (.in_A(in_A[67]), .in_B(in_B[67]), .in_CI(nC67), .out_S(out_S[67]), .out_CO(nC68));
  VFA U68 (.in_A(in_A[68]), .in_B(in_B[68]), .in_CI(nC68), .out_S(out_S[68]), .out_CO(nC69));
  VFA U69 (.in_A(in_A[69]), .in_B(in_B[69]), .in_CI(nC69), .out_S(out_S[69]), .out_CO(nC70));
  VFA U70 (.in_A(in_A[70]), .in_B(in_B[70]), .in_CI(nC70), .out_S(out_S[70]), .out_CO(nC71));
  VFA U71 (.in_A(in_A[71]), .in_B(in_B[71]), .in_CI(nC71), .out_S(out_S[71]), .out_CO(nC72));
  VFA U72 (.in_A(in_A[72]), .in_B(in_B[72]), .in_CI(nC72), .out_S(out_S[72]), .out_CO(nC73));
  VFA U73 (.in_A(in_A[73]), .in_B(in_B[73]), .in_CI(nC73), .out_S(out_S[73]), .out_CO(nC74));
  VFA U74 (.in_A(in_A[74]), .in_B(in_B[74]), .in_CI(nC74), .out_S(out_S[74]), .out_CO(nC75));
  VFA U75 (.in_A(in_A[75]), .in_B(in_B[75]), .in_CI(nC75), .out_S(out_S[75]), .out_CO(nC76));
  VFA U76 (.in_A(in_A[76]), .in_B(in_B[76]), .in_CI(nC76), .out_S(out_S[76]), .out_CO(nC77));
  VFA U77 (.in_A(in_A[77]), .in_B(in_B[77]), .in_CI(nC77), .out_S(out_S[77]), .out_CO(nC78));
  VFA U78 (.in_A(in_A[78]), .in_B(in_B[78]), .in_CI(nC78), .out_S(out_S[78]), .out_CO(nC79));
  VFA U79 (.in_A(in_A[79]), .in_B(in_B[79]), .in_CI(nC79), .out_S(out_S[79]), .out_CO(nC80));
  VFA U80 (.in_A(in_A[80]), .in_B(in_B[80]), .in_CI(nC80), .out_S(out_S[80]), .out_CO(nC81));
  VFA U81 (.in_A(in_A[81]), .in_B(in_B[81]), .in_CI(nC81), .out_S(out_S[81]), .out_CO(nC82));
  VFA U82 (.in_A(in_A[82]), .in_B(in_B[82]), .in_CI(nC82), .out_S(out_S[82]), .out_CO(nC83));
  VFA U83 (.in_A(in_A[83]), .in_B(in_B[83]), .in_CI(nC83), .out_S(out_S[83]), .out_CO(nC84));
  VFA U84 (.in_A(in_A[84]), .in_B(in_B[84]), .in_CI(nC84), .out_S(out_S[84]), .out_CO(nC85));
  VFA U85 (.in_A(in_A[85]), .in_B(in_B[85]), .in_CI(nC85), .out_S(out_S[85]), .out_CO(nC86));
  VFA U86 (.in_A(in_A[86]), .in_B(in_B[86]), .in_CI(nC86), .out_S(out_S[86]), .out_CO(nC87));
  VFA U87 (.in_A(in_A[87]), .in_B(in_B[87]), .in_CI(nC87), .out_S(out_S[87]), .out_CO(nC88));
  VFA U88 (.in_A(in_A[88]), .in_B(in_B[88]), .in_CI(nC88), .out_S(out_S[88]), .out_CO(nC89));
  VFA U89 (.in_A(in_A[89]), .in_B(in_B[89]), .in_CI(nC89), .out_S(out_S[89]), .out_CO(nC90));
  VFA U90 (.in_A(in_A[90]), .in_B(in_B[90]), .in_CI(nC90), .out_S(out_S[90]), .out_CO(nC91));
  VFA U91 (.in_A(in_A[91]), .in_B(in_B[91]), .in_CI(nC91), .out_S(out_S[91]), .out_CO(nC92));
  VFA U92 (.in_A(in_A[92]), .in_B(in_B[92]), .in_CI(nC92), .out_S(out_S[92]), .out_CO(nC93));
  VFA U93 (.in_A(in_A[93]), .in_B(in_B[93]), .in_CI(nC93), .out_S(out_S[93]), .out_CO(nC94));
  VFA U94 (.in_A(in_A[94]), .in_B(in_B[94]), .in_CI(nC94), .out_S(out_S[94]), .out_CO(nC95));
  VFA U95 (.in_A(in_A[95]), .in_B(in_B[95]), .in_CI(nC95), .out_S(out_S[95]), .out_CO(nC96));
  VFA U96 (.in_A(in_A[96]), .in_B(in_B[96]), .in_CI(nC96), .out_S(out_S[96]), .out_CO(nC97));
  VFA U97 (.in_A(in_A[97]), .in_B(in_B[97]), .in_CI(nC97), .out_S(out_S[97]), .out_CO(nC98));
  VFA U98 (.in_A(in_A[98]), .in_B(in_B[98]), .in_CI(nC98), .out_S(out_S[98]), .out_CO(nC99));
  VFA U99 (.in_A(in_A[99]), .in_B(in_B[99]), .in_CI(nC99), .out_S(out_S[99]), .out_CO(nC100));
  VFA U100 (.in_A(in_A[100]), .in_B(in_B[100]), .in_CI(nC100), .out_S(out_S[100]), .out_CO(nC101));
  VFA U101 (.in_A(in_A[101]), .in_B(in_B[101]), .in_CI(nC101), .out_S(out_S[101]), .out_CO(nC102));
  VFA U102 (.in_A(in_A[102]), .in_B(in_B[102]), .in_CI(nC102), .out_S(out_S[102]), .out_CO(nC103));
  VFA U103 (.in_A(in_A[103]), .in_B(in_B[103]), .in_CI(nC103), .out_S(out_S[103]), .out_CO(nC104));
  VFA U104 (.in_A(in_A[104]), .in_B(in_B[104]), .in_CI(nC104), .out_S(out_S[104]), .out_CO(nC105));
  VFA U105 (.in_A(in_A[105]), .in_B(in_B[105]), .in_CI(nC105), .out_S(out_S[105]), .out_CO(nC106));
  VFA U106 (.in_A(in_A[106]), .in_B(in_B[106]), .in_CI(nC106), .out_S(out_S[106]), .out_CO(nC107));
  VFA U107 (.in_A(in_A[107]), .in_B(in_B[107]), .in_CI(nC107), .out_S(out_S[107]), .out_CO(nC108));
  VFA U108 (.in_A(in_A[108]), .in_B(in_B[108]), .in_CI(nC108), .out_S(out_S[108]), .out_CO(nC109));
  VFA U109 (.in_A(in_A[109]), .in_B(in_B[109]), .in_CI(nC109), .out_S(out_S[109]), .out_CO(nC110));
  VFA U110 (.in_A(in_A[110]), .in_B(in_B[110]), .in_CI(nC110), .out_S(out_S[110]), .out_CO(nC111));
  VFA U111 (.in_A(in_A[111]), .in_B(in_B[111]), .in_CI(nC111), .out_S(out_S[111]), .out_CO(nC112));
  VFA U112 (.in_A(in_A[112]), .in_B(in_B[112]), .in_CI(nC112), .out_S(out_S[112]), .out_CO(nC113));
  VFA U113 (.in_A(in_A[113]), .in_B(in_B[113]), .in_CI(nC113), .out_S(out_S[113]), .out_CO(nC114));
  VFA U114 (.in_A(in_A[114]), .in_B(in_B[114]), .in_CI(nC114), .out_S(out_S[114]), .out_CO(nC115));
  VFA U115 (.in_A(in_A[115]), .in_B(in_B[115]), .in_CI(nC115), .out_S(out_S[115]), .out_CO(nC116));
  VFA U116 (.in_A(in_A[116]), .in_B(in_B[116]), .in_CI(nC116), .out_S(out_S[116]), .out_CO(nC117));
  VFA U117 (.in_A(in_A[117]), .in_B(in_B[117]), .in_CI(nC117), .out_S(out_S[117]), .out_CO(nC118));
  VFA U118 (.in_A(in_A[118]), .in_B(in_B[118]), .in_CI(nC118), .out_S(out_S[118]), .out_CO(nC119));
  VFA U119 (.in_A(in_A[119]), .in_B(in_B[119]), .in_CI(nC119), .out_S(out_S[119]), .out_CO(nC120));
  VFA U120 (.in_A(in_A[120]), .in_B(in_B[120]), .in_CI(nC120), .out_S(out_S[120]), .out_CO(nC121));
  VFA U121 (.in_A(in_A[121]), .in_B(in_B[121]), .in_CI(nC121), .out_S(out_S[121]), .out_CO(nC122));
  VFA U122 (.in_A(in_A[122]), .in_B(in_B[122]), .in_CI(nC122), .out_S(out_S[122]), .out_CO(nC123));
  VFA U123 (.in_A(in_A[123]), .in_B(in_B[123]), .in_CI(nC123), .out_S(out_S[123]), .out_CO(nC124));
  VFA U124 (.in_A(in_A[124]), .in_B(in_B[124]), .in_CI(nC124), .out_S(out_S[124]), .out_CO(nC125));
  VFA U125 (.in_A(in_A[125]), .in_B(in_B[125]), .in_CI(nC125), .out_S(out_S[125]), .out_CO(nC126));
  VFA U126 (.in_A(in_A[126]), .in_B(in_B[126]), .in_CI(nC126), .out_S(out_S[126]), .out_CO(nC127));
  VFA U127 (.in_A(in_A[127]), .in_B(in_B[127]), .in_CI(nC127), .out_S(out_S[127]), .out_CO(nC128));
  VFA U128 (.in_A(in_A[128]), .in_B(in_B[128]), .in_CI(nC128), .out_S(out_S[128]), .out_CO(nC129));
  VFA U129 (.in_A(in_A[129]), .in_B(in_B[129]), .in_CI(nC129), .out_S(out_S[129]), .out_CO(nC130));
  VFA U130 (.in_A(in_A[130]), .in_B(in_B[130]), .in_CI(nC130), .out_S(out_S[130]), .out_CO(nC131));
  VFA U131 (.in_A(in_A[131]), .in_B(in_B[131]), .in_CI(nC131), .out_S(out_S[131]), .out_CO(nC132));
  VFA U132 (.in_A(in_A[132]), .in_B(in_B[132]), .in_CI(nC132), .out_S(out_S[132]), .out_CO(nC133));
  VFA U133 (.in_A(in_A[133]), .in_B(in_B[133]), .in_CI(nC133), .out_S(out_S[133]), .out_CO(nC134));
  VFA U134 (.in_A(in_A[134]), .in_B(in_B[134]), .in_CI(nC134), .out_S(out_S[134]), .out_CO(nC135));
  VFA U135 (.in_A(in_A[135]), .in_B(in_B[135]), .in_CI(nC135), .out_S(out_S[135]), .out_CO(nC136));
  VFA U136 (.in_A(in_A[136]), .in_B(in_B[136]), .in_CI(nC136), .out_S(out_S[136]), .out_CO(nC137));
  VFA U137 (.in_A(in_A[137]), .in_B(in_B[137]), .in_CI(nC137), .out_S(out_S[137]), .out_CO(nC138));
  VFA U138 (.in_A(in_A[138]), .in_B(in_B[138]), .in_CI(nC138), .out_S(out_S[138]), .out_CO(nC139));
  VFA U139 (.in_A(in_A[139]), .in_B(in_B[139]), .in_CI(nC139), .out_S(out_S[139]), .out_CO(nC140));
  VFA U140 (.in_A(in_A[140]), .in_B(in_B[140]), .in_CI(nC140), .out_S(out_S[140]), .out_CO(nC141));
  VFA U141 (.in_A(in_A[141]), .in_B(in_B[141]), .in_CI(nC141), .out_S(out_S[141]), .out_CO(nC142));
  VFA U142 (.in_A(in_A[142]), .in_B(in_B[142]), .in_CI(nC142), .out_S(out_S[142]), .out_CO(nC143));
  VFA U143 (.in_A(in_A[143]), .in_B(in_B[143]), .in_CI(nC143), .out_S(out_S[143]), .out_CO(nC144));
  VFA U144 (.in_A(in_A[144]), .in_B(in_B[144]), .in_CI(nC144), .out_S(out_S[144]), .out_CO(nC145));
  VFA U145 (.in_A(in_A[145]), .in_B(in_B[145]), .in_CI(nC145), .out_S(out_S[145]), .out_CO(nC146));
  VFA U146 (.in_A(in_A[146]), .in_B(in_B[146]), .in_CI(nC146), .out_S(out_S[146]), .out_CO(nC147));
  VFA U147 (.in_A(in_A[147]), .in_B(in_B[147]), .in_CI(nC147), .out_S(out_S[147]), .out_CO(nC148));
  VFA U148 (.in_A(in_A[148]), .in_B(in_B[148]), .in_CI(nC148), .out_S(out_S[148]), .out_CO(nC149));
  VFA U149 (.in_A(in_A[149]), .in_B(in_B[149]), .in_CI(nC149), .out_S(out_S[149]), .out_CO(nC150));
  VFA U150 (.in_A(in_A[150]), .in_B(in_B[150]), .in_CI(nC150), .out_S(out_S[150]), .out_CO(nC151));
  VFA U151 (.in_A(in_A[151]), .in_B(in_B[151]), .in_CI(nC151), .out_S(out_S[151]), .out_CO(nC152));
  VFA U152 (.in_A(in_A[152]), .in_B(in_B[152]), .in_CI(nC152), .out_S(out_S[152]), .out_CO(nC153));
  VFA U153 (.in_A(in_A[153]), .in_B(in_B[153]), .in_CI(nC153), .out_S(out_S[153]), .out_CO(nC154));
  VFA U154 (.in_A(in_A[154]), .in_B(in_B[154]), .in_CI(nC154), .out_S(out_S[154]), .out_CO(nC155));
  VFA U155 (.in_A(in_A[155]), .in_B(in_B[155]), .in_CI(nC155), .out_S(out_S[155]), .out_CO(nC156));
  VFA U156 (.in_A(in_A[156]), .in_B(in_B[156]), .in_CI(nC156), .out_S(out_S[156]), .out_CO(nC157));
  VFA U157 (.in_A(in_A[157]), .in_B(in_B[157]), .in_CI(nC157), .out_S(out_S[157]), .out_CO(nC158));
  VFA U158 (.in_A(in_A[158]), .in_B(in_B[158]), .in_CI(nC158), .out_S(out_S[158]), .out_CO(nC159));
  VFA U159 (.in_A(in_A[159]), .in_B(in_B[159]), .in_CI(nC159), .out_S(out_S[159]), .out_CO(nC160));
  VFA U160 (.in_A(in_A[160]), .in_B(in_B[160]), .in_CI(nC160), .out_S(out_S[160]), .out_CO(nC161));
  VFA U161 (.in_A(in_A[161]), .in_B(in_B[161]), .in_CI(nC161), .out_S(out_S[161]), .out_CO(nC162));
  VFA U162 (.in_A(in_A[162]), .in_B(in_B[162]), .in_CI(nC162), .out_S(out_S[162]), .out_CO(nC163));
  VFA U163 (.in_A(in_A[163]), .in_B(in_B[163]), .in_CI(nC163), .out_S(out_S[163]), .out_CO(nC164));
  VFA U164 (.in_A(in_A[164]), .in_B(in_B[164]), .in_CI(nC164), .out_S(out_S[164]), .out_CO(nC165));
  VFA U165 (.in_A(in_A[165]), .in_B(in_B[165]), .in_CI(nC165), .out_S(out_S[165]), .out_CO(nC166));
  VFA U166 (.in_A(in_A[166]), .in_B(in_B[166]), .in_CI(nC166), .out_S(out_S[166]), .out_CO(nC167));
  VFA U167 (.in_A(in_A[167]), .in_B(in_B[167]), .in_CI(nC167), .out_S(out_S[167]), .out_CO(nC168));
  VFA U168 (.in_A(in_A[168]), .in_B(in_B[168]), .in_CI(nC168), .out_S(out_S[168]), .out_CO(nC169));
  VFA U169 (.in_A(in_A[169]), .in_B(in_B[169]), .in_CI(nC169), .out_S(out_S[169]), .out_CO(nC170));
  VFA U170 (.in_A(in_A[170]), .in_B(in_B[170]), .in_CI(nC170), .out_S(out_S[170]), .out_CO(nC171));
  VFA U171 (.in_A(in_A[171]), .in_B(in_B[171]), .in_CI(nC171), .out_S(out_S[171]), .out_CO(nC172));
  VFA U172 (.in_A(in_A[172]), .in_B(in_B[172]), .in_CI(nC172), .out_S(out_S[172]), .out_CO(nC173));
  VFA U173 (.in_A(in_A[173]), .in_B(in_B[173]), .in_CI(nC173), .out_S(out_S[173]), .out_CO(nC174));
  VFA U174 (.in_A(in_A[174]), .in_B(in_B[174]), .in_CI(nC174), .out_S(out_S[174]), .out_CO(nC175));
  VFA U175 (.in_A(in_A[175]), .in_B(in_B[175]), .in_CI(nC175), .out_S(out_S[175]), .out_CO(nC176));
  VFA U176 (.in_A(in_A[176]), .in_B(in_B[176]), .in_CI(nC176), .out_S(out_S[176]), .out_CO(nC177));
  VFA U177 (.in_A(in_A[177]), .in_B(in_B[177]), .in_CI(nC177), .out_S(out_S[177]), .out_CO(nC178));
  VFA U178 (.in_A(in_A[178]), .in_B(in_B[178]), .in_CI(nC178), .out_S(out_S[178]), .out_CO(nC179));
  VFA U179 (.in_A(in_A[179]), .in_B(in_B[179]), .in_CI(nC179), .out_S(out_S[179]), .out_CO(nC180));
  VFA U180 (.in_A(in_A[180]), .in_B(in_B[180]), .in_CI(nC180), .out_S(out_S[180]), .out_CO(nC181));
  VFA U181 (.in_A(in_A[181]), .in_B(in_B[181]), .in_CI(nC181), .out_S(out_S[181]), .out_CO(nC182));
  VFA U182 (.in_A(in_A[182]), .in_B(in_B[182]), .in_CI(nC182), .out_S(out_S[182]), .out_CO(nC183));
  VFA U183 (.in_A(in_A[183]), .in_B(in_B[183]), .in_CI(nC183), .out_S(out_S[183]), .out_CO(nC184));
  VFA U184 (.in_A(in_A[184]), .in_B(in_B[184]), .in_CI(nC184), .out_S(out_S[184]), .out_CO(nC185));
  VFA U185 (.in_A(in_A[185]), .in_B(in_B[185]), .in_CI(nC185), .out_S(out_S[185]), .out_CO(nC186));
  VFA U186 (.in_A(in_A[186]), .in_B(in_B[186]), .in_CI(nC186), .out_S(out_S[186]), .out_CO(nC187));
  VFA U187 (.in_A(in_A[187]), .in_B(in_B[187]), .in_CI(nC187), .out_S(out_S[187]), .out_CO(nC188));
  VFA U188 (.in_A(in_A[188]), .in_B(in_B[188]), .in_CI(nC188), .out_S(out_S[188]), .out_CO(nC189));
  VFA U189 (.in_A(in_A[189]), .in_B(in_B[189]), .in_CI(nC189), .out_S(out_S[189]), .out_CO(nC190));
  VFA U190 (.in_A(in_A[190]), .in_B(in_B[190]), .in_CI(nC190), .out_S(out_S[190]), .out_CO(nC191));
  VFA U191 (.in_A(in_A[191]), .in_B(in_B[191]), .in_CI(nC191), .out_S(out_S[191]), .out_CO(nC192));
  VFA U192 (.in_A(in_A[192]), .in_B(in_B[192]), .in_CI(nC192), .out_S(out_S[192]), .out_CO(nC193));
  VFA U193 (.in_A(in_A[193]), .in_B(in_B[193]), .in_CI(nC193), .out_S(out_S[193]), .out_CO(nC194));
  VFA U194 (.in_A(in_A[194]), .in_B(in_B[194]), .in_CI(nC194), .out_S(out_S[194]), .out_CO(nC195));
  VFA U195 (.in_A(in_A[195]), .in_B(in_B[195]), .in_CI(nC195), .out_S(out_S[195]), .out_CO(nC196));
  VFA U196 (.in_A(in_A[196]), .in_B(in_B[196]), .in_CI(nC196), .out_S(out_S[196]), .out_CO(nC197));
  VFA U197 (.in_A(in_A[197]), .in_B(in_B[197]), .in_CI(nC197), .out_S(out_S[197]), .out_CO(nC198));
  VFA U198 (.in_A(in_A[198]), .in_B(in_B[198]), .in_CI(nC198), .out_S(out_S[198]), .out_CO(nC199));
  VFA U199 (.in_A(in_A[199]), .in_B(in_B[199]), .in_CI(nC199), .out_S(out_S[199]), .out_CO(nC200));
  VFA U200 (.in_A(in_A[200]), .in_B(in_B[200]), .in_CI(nC200), .out_S(out_S[200]), .out_CO(nC201));
  VFA U201 (.in_A(in_A[201]), .in_B(in_B[201]), .in_CI(nC201), .out_S(out_S[201]), .out_CO(nC202));
  VFA U202 (.in_A(in_A[202]), .in_B(in_B[202]), .in_CI(nC202), .out_S(out_S[202]), .out_CO(nC203));
  VFA U203 (.in_A(in_A[203]), .in_B(in_B[203]), .in_CI(nC203), .out_S(out_S[203]), .out_CO(nC204));
  VFA U204 (.in_A(in_A[204]), .in_B(in_B[204]), .in_CI(nC204), .out_S(out_S[204]), .out_CO(nC205));
  VFA U205 (.in_A(in_A[205]), .in_B(in_B[205]), .in_CI(nC205), .out_S(out_S[205]), .out_CO(nC206));
  VFA U206 (.in_A(in_A[206]), .in_B(in_B[206]), .in_CI(nC206), .out_S(out_S[206]), .out_CO(nC207));
  VFA U207 (.in_A(in_A[207]), .in_B(in_B[207]), .in_CI(nC207), .out_S(out_S[207]), .out_CO(nC208));
  VFA U208 (.in_A(in_A[208]), .in_B(in_B[208]), .in_CI(nC208), .out_S(out_S[208]), .out_CO(nC209));
  VFA U209 (.in_A(in_A[209]), .in_B(in_B[209]), .in_CI(nC209), .out_S(out_S[209]), .out_CO(nC210));
  VFA U210 (.in_A(in_A[210]), .in_B(in_B[210]), .in_CI(nC210), .out_S(out_S[210]), .out_CO(nC211));
  VFA U211 (.in_A(in_A[211]), .in_B(in_B[211]), .in_CI(nC211), .out_S(out_S[211]), .out_CO(nC212));
  VFA U212 (.in_A(in_A[212]), .in_B(in_B[212]), .in_CI(nC212), .out_S(out_S[212]), .out_CO(nC213));
  VFA U213 (.in_A(in_A[213]), .in_B(in_B[213]), .in_CI(nC213), .out_S(out_S[213]), .out_CO(nC214));
  VFA U214 (.in_A(in_A[214]), .in_B(in_B[214]), .in_CI(nC214), .out_S(out_S[214]), .out_CO(nC215));
  VFA U215 (.in_A(in_A[215]), .in_B(in_B[215]), .in_CI(nC215), .out_S(out_S[215]), .out_CO(nC216));
  VFA U216 (.in_A(in_A[216]), .in_B(in_B[216]), .in_CI(nC216), .out_S(out_S[216]), .out_CO(nC217));
  VFA U217 (.in_A(in_A[217]), .in_B(in_B[217]), .in_CI(nC217), .out_S(out_S[217]), .out_CO(nC218));
  VFA U218 (.in_A(in_A[218]), .in_B(in_B[218]), .in_CI(nC218), .out_S(out_S[218]), .out_CO(nC219));
  VFA U219 (.in_A(in_A[219]), .in_B(in_B[219]), .in_CI(nC219), .out_S(out_S[219]), .out_CO(nC220));
  VFA U220 (.in_A(in_A[220]), .in_B(in_B[220]), .in_CI(nC220), .out_S(out_S[220]), .out_CO(nC221));
  VFA U221 (.in_A(in_A[221]), .in_B(in_B[221]), .in_CI(nC221), .out_S(out_S[221]), .out_CO(nC222));
  VFA U222 (.in_A(in_A[222]), .in_B(in_B[222]), .in_CI(nC222), .out_S(out_S[222]), .out_CO(nC223));
  VFA U223 (.in_A(in_A[223]), .in_B(in_B[223]), .in_CI(nC223), .out_S(out_S[223]), .out_CO(nC224));
  VFA U224 (.in_A(in_A[224]), .in_B(in_B[224]), .in_CI(nC224), .out_S(out_S[224]), .out_CO(nC225));
  VFA U225 (.in_A(in_A[225]), .in_B(in_B[225]), .in_CI(nC225), .out_S(out_S[225]), .out_CO(nC226));
  VFA U226 (.in_A(in_A[226]), .in_B(in_B[226]), .in_CI(nC226), .out_S(out_S[226]), .out_CO(nC227));
  VFA U227 (.in_A(in_A[227]), .in_B(in_B[227]), .in_CI(nC227), .out_S(out_S[227]), .out_CO(nC228));
  VFA U228 (.in_A(in_A[228]), .in_B(in_B[228]), .in_CI(nC228), .out_S(out_S[228]), .out_CO(nC229));
  VFA U229 (.in_A(in_A[229]), .in_B(in_B[229]), .in_CI(nC229), .out_S(out_S[229]), .out_CO(nC230));
  VFA U230 (.in_A(in_A[230]), .in_B(in_B[230]), .in_CI(nC230), .out_S(out_S[230]), .out_CO(nC231));
  VFA U231 (.in_A(in_A[231]), .in_B(in_B[231]), .in_CI(nC231), .out_S(out_S[231]), .out_CO(nC232));
  VFA U232 (.in_A(in_A[232]), .in_B(in_B[232]), .in_CI(nC232), .out_S(out_S[232]), .out_CO(nC233));
  VFA U233 (.in_A(in_A[233]), .in_B(in_B[233]), .in_CI(nC233), .out_S(out_S[233]), .out_CO(nC234));
  VFA U234 (.in_A(in_A[234]), .in_B(in_B[234]), .in_CI(nC234), .out_S(out_S[234]), .out_CO(nC235));
  VFA U235 (.in_A(in_A[235]), .in_B(in_B[235]), .in_CI(nC235), .out_S(out_S[235]), .out_CO(nC236));
  VFA U236 (.in_A(in_A[236]), .in_B(in_B[236]), .in_CI(nC236), .out_S(out_S[236]), .out_CO(nC237));
  VFA U237 (.in_A(in_A[237]), .in_B(in_B[237]), .in_CI(nC237), .out_S(out_S[237]), .out_CO(nC238));
  VFA U238 (.in_A(in_A[238]), .in_B(in_B[238]), .in_CI(nC238), .out_S(out_S[238]), .out_CO(nC239));
  VFA U239 (.in_A(in_A[239]), .in_B(in_B[239]), .in_CI(nC239), .out_S(out_S[239]), .out_CO(nC240));
  VFA U240 (.in_A(in_A[240]), .in_B(in_B[240]), .in_CI(nC240), .out_S(out_S[240]), .out_CO(nC241));
  VFA U241 (.in_A(in_A[241]), .in_B(in_B[241]), .in_CI(nC241), .out_S(out_S[241]), .out_CO(nC242));
  VFA U242 (.in_A(in_A[242]), .in_B(in_B[242]), .in_CI(nC242), .out_S(out_S[242]), .out_CO(nC243));
  VFA U243 (.in_A(in_A[243]), .in_B(in_B[243]), .in_CI(nC243), .out_S(out_S[243]), .out_CO(nC244));
  VFA U244 (.in_A(in_A[244]), .in_B(in_B[244]), .in_CI(nC244), .out_S(out_S[244]), .out_CO(nC245));
  VFA U245 (.in_A(in_A[245]), .in_B(in_B[245]), .in_CI(nC245), .out_S(out_S[245]), .out_CO(nC246));
  VFA U246 (.in_A(in_A[246]), .in_B(in_B[246]), .in_CI(nC246), .out_S(out_S[246]), .out_CO(nC247));
  VFA U247 (.in_A(in_A[247]), .in_B(in_B[247]), .in_CI(nC247), .out_S(out_S[247]), .out_CO(nC248));
  VFA U248 (.in_A(in_A[248]), .in_B(in_B[248]), .in_CI(nC248), .out_S(out_S[248]), .out_CO(nC249));
  VFA U249 (.in_A(in_A[249]), .in_B(in_B[249]), .in_CI(nC249), .out_S(out_S[249]), .out_CO(nC250));
  VFA U250 (.in_A(in_A[250]), .in_B(in_B[250]), .in_CI(nC250), .out_S(out_S[250]), .out_CO(nC251));
  VFA U251 (.in_A(in_A[251]), .in_B(in_B[251]), .in_CI(nC251), .out_S(out_S[251]), .out_CO(nC252));
  VFA U252 (.in_A(in_A[252]), .in_B(in_B[252]), .in_CI(nC252), .out_S(out_S[252]), .out_CO(nC253));
  VFA U253 (.in_A(in_A[253]), .in_B(in_B[253]), .in_CI(nC253), .out_S(out_S[253]), .out_CO(nC254));
  VFA U254 (.in_A(in_A[254]), .in_B(in_B[254]), .in_CI(nC254), .out_S(out_S[254]), .out_CO(nC255));
  VFA U255 (.in_A(in_A[255]), .in_B(in_B[255]), .in_CI(nC255), .out_S(out_S[255]), .out_CO(out_CO));
endmodule

