module VFA (in_A, in_B, in_CI, out_S, out_CO);
  input in_A, in_B, in_CI;
  output out_S, out_CO;

  assign out_S = in_A ^ in_B ^ in_CI;
  assign out_CO = (in_A & in_B) | (in_B & in_CI) | (in_CI & in_A);
endmodule



module VRCA_128 (in_A, in_B, in_CI, out_S, out_CO);
  input [127:0] in_A, in_B;
  input in_CI;
  output [127:0] out_S;
  output out_CO;

  VFA U0 (.in_A(in_A[0]), .in_B(in_B[0]), .in_CI(in_CI), .out_S(out_S[0]), .out_CO(nC1));
  VFA U1 (.in_A(in_A[1]), .in_B(in_B[1]), .in_CI(nC1), .out_S(out_S[1]), .out_CO(nC2));
  VFA U2 (.in_A(in_A[2]), .in_B(in_B[2]), .in_CI(nC2), .out_S(out_S[2]), .out_CO(nC3));
  VFA U3 (.in_A(in_A[3]), .in_B(in_B[3]), .in_CI(nC3), .out_S(out_S[3]), .out_CO(nC4));
  VFA U4 (.in_A(in_A[4]), .in_B(in_B[4]), .in_CI(nC4), .out_S(out_S[4]), .out_CO(nC5));
  VFA U5 (.in_A(in_A[5]), .in_B(in_B[5]), .in_CI(nC5), .out_S(out_S[5]), .out_CO(nC6));
  VFA U6 (.in_A(in_A[6]), .in_B(in_B[6]), .in_CI(nC6), .out_S(out_S[6]), .out_CO(nC7));
  VFA U7 (.in_A(in_A[7]), .in_B(in_B[7]), .in_CI(nC7), .out_S(out_S[7]), .out_CO(nC8));
  VFA U8 (.in_A(in_A[8]), .in_B(in_B[8]), .in_CI(nC8), .out_S(out_S[8]), .out_CO(nC9));
  VFA U9 (.in_A(in_A[9]), .in_B(in_B[9]), .in_CI(nC9), .out_S(out_S[9]), .out_CO(nC10));
  VFA U10 (.in_A(in_A[10]), .in_B(in_B[10]), .in_CI(nC10), .out_S(out_S[10]), .out_CO(nC11));
  VFA U11 (.in_A(in_A[11]), .in_B(in_B[11]), .in_CI(nC11), .out_S(out_S[11]), .out_CO(nC12));
  VFA U12 (.in_A(in_A[12]), .in_B(in_B[12]), .in_CI(nC12), .out_S(out_S[12]), .out_CO(nC13));
  VFA U13 (.in_A(in_A[13]), .in_B(in_B[13]), .in_CI(nC13), .out_S(out_S[13]), .out_CO(nC14));
  VFA U14 (.in_A(in_A[14]), .in_B(in_B[14]), .in_CI(nC14), .out_S(out_S[14]), .out_CO(nC15));
  VFA U15 (.in_A(in_A[15]), .in_B(in_B[15]), .in_CI(nC15), .out_S(out_S[15]), .out_CO(nC16));
  VFA U16 (.in_A(in_A[16]), .in_B(in_B[16]), .in_CI(nC16), .out_S(out_S[16]), .out_CO(nC17));
  VFA U17 (.in_A(in_A[17]), .in_B(in_B[17]), .in_CI(nC17), .out_S(out_S[17]), .out_CO(nC18));
  VFA U18 (.in_A(in_A[18]), .in_B(in_B[18]), .in_CI(nC18), .out_S(out_S[18]), .out_CO(nC19));
  VFA U19 (.in_A(in_A[19]), .in_B(in_B[19]), .in_CI(nC19), .out_S(out_S[19]), .out_CO(nC20));
  VFA U20 (.in_A(in_A[20]), .in_B(in_B[20]), .in_CI(nC20), .out_S(out_S[20]), .out_CO(nC21));
  VFA U21 (.in_A(in_A[21]), .in_B(in_B[21]), .in_CI(nC21), .out_S(out_S[21]), .out_CO(nC22));
  VFA U22 (.in_A(in_A[22]), .in_B(in_B[22]), .in_CI(nC22), .out_S(out_S[22]), .out_CO(nC23));
  VFA U23 (.in_A(in_A[23]), .in_B(in_B[23]), .in_CI(nC23), .out_S(out_S[23]), .out_CO(nC24));
  VFA U24 (.in_A(in_A[24]), .in_B(in_B[24]), .in_CI(nC24), .out_S(out_S[24]), .out_CO(nC25));
  VFA U25 (.in_A(in_A[25]), .in_B(in_B[25]), .in_CI(nC25), .out_S(out_S[25]), .out_CO(nC26));
  VFA U26 (.in_A(in_A[26]), .in_B(in_B[26]), .in_CI(nC26), .out_S(out_S[26]), .out_CO(nC27));
  VFA U27 (.in_A(in_A[27]), .in_B(in_B[27]), .in_CI(nC27), .out_S(out_S[27]), .out_CO(nC28));
  VFA U28 (.in_A(in_A[28]), .in_B(in_B[28]), .in_CI(nC28), .out_S(out_S[28]), .out_CO(nC29));
  VFA U29 (.in_A(in_A[29]), .in_B(in_B[29]), .in_CI(nC29), .out_S(out_S[29]), .out_CO(nC30));
  VFA U30 (.in_A(in_A[30]), .in_B(in_B[30]), .in_CI(nC30), .out_S(out_S[30]), .out_CO(nC31));
  VFA U31 (.in_A(in_A[31]), .in_B(in_B[31]), .in_CI(nC31), .out_S(out_S[31]), .out_CO(nC32));
  VFA U32 (.in_A(in_A[32]), .in_B(in_B[32]), .in_CI(nC32), .out_S(out_S[32]), .out_CO(nC33));
  VFA U33 (.in_A(in_A[33]), .in_B(in_B[33]), .in_CI(nC33), .out_S(out_S[33]), .out_CO(nC34));
  VFA U34 (.in_A(in_A[34]), .in_B(in_B[34]), .in_CI(nC34), .out_S(out_S[34]), .out_CO(nC35));
  VFA U35 (.in_A(in_A[35]), .in_B(in_B[35]), .in_CI(nC35), .out_S(out_S[35]), .out_CO(nC36));
  VFA U36 (.in_A(in_A[36]), .in_B(in_B[36]), .in_CI(nC36), .out_S(out_S[36]), .out_CO(nC37));
  VFA U37 (.in_A(in_A[37]), .in_B(in_B[37]), .in_CI(nC37), .out_S(out_S[37]), .out_CO(nC38));
  VFA U38 (.in_A(in_A[38]), .in_B(in_B[38]), .in_CI(nC38), .out_S(out_S[38]), .out_CO(nC39));
  VFA U39 (.in_A(in_A[39]), .in_B(in_B[39]), .in_CI(nC39), .out_S(out_S[39]), .out_CO(nC40));
  VFA U40 (.in_A(in_A[40]), .in_B(in_B[40]), .in_CI(nC40), .out_S(out_S[40]), .out_CO(nC41));
  VFA U41 (.in_A(in_A[41]), .in_B(in_B[41]), .in_CI(nC41), .out_S(out_S[41]), .out_CO(nC42));
  VFA U42 (.in_A(in_A[42]), .in_B(in_B[42]), .in_CI(nC42), .out_S(out_S[42]), .out_CO(nC43));
  VFA U43 (.in_A(in_A[43]), .in_B(in_B[43]), .in_CI(nC43), .out_S(out_S[43]), .out_CO(nC44));
  VFA U44 (.in_A(in_A[44]), .in_B(in_B[44]), .in_CI(nC44), .out_S(out_S[44]), .out_CO(nC45));
  VFA U45 (.in_A(in_A[45]), .in_B(in_B[45]), .in_CI(nC45), .out_S(out_S[45]), .out_CO(nC46));
  VFA U46 (.in_A(in_A[46]), .in_B(in_B[46]), .in_CI(nC46), .out_S(out_S[46]), .out_CO(nC47));
  VFA U47 (.in_A(in_A[47]), .in_B(in_B[47]), .in_CI(nC47), .out_S(out_S[47]), .out_CO(nC48));
  VFA U48 (.in_A(in_A[48]), .in_B(in_B[48]), .in_CI(nC48), .out_S(out_S[48]), .out_CO(nC49));
  VFA U49 (.in_A(in_A[49]), .in_B(in_B[49]), .in_CI(nC49), .out_S(out_S[49]), .out_CO(nC50));
  VFA U50 (.in_A(in_A[50]), .in_B(in_B[50]), .in_CI(nC50), .out_S(out_S[50]), .out_CO(nC51));
  VFA U51 (.in_A(in_A[51]), .in_B(in_B[51]), .in_CI(nC51), .out_S(out_S[51]), .out_CO(nC52));
  VFA U52 (.in_A(in_A[52]), .in_B(in_B[52]), .in_CI(nC52), .out_S(out_S[52]), .out_CO(nC53));
  VFA U53 (.in_A(in_A[53]), .in_B(in_B[53]), .in_CI(nC53), .out_S(out_S[53]), .out_CO(nC54));
  VFA U54 (.in_A(in_A[54]), .in_B(in_B[54]), .in_CI(nC54), .out_S(out_S[54]), .out_CO(nC55));
  VFA U55 (.in_A(in_A[55]), .in_B(in_B[55]), .in_CI(nC55), .out_S(out_S[55]), .out_CO(nC56));
  VFA U56 (.in_A(in_A[56]), .in_B(in_B[56]), .in_CI(nC56), .out_S(out_S[56]), .out_CO(nC57));
  VFA U57 (.in_A(in_A[57]), .in_B(in_B[57]), .in_CI(nC57), .out_S(out_S[57]), .out_CO(nC58));
  VFA U58 (.in_A(in_A[58]), .in_B(in_B[58]), .in_CI(nC58), .out_S(out_S[58]), .out_CO(nC59));
  VFA U59 (.in_A(in_A[59]), .in_B(in_B[59]), .in_CI(nC59), .out_S(out_S[59]), .out_CO(nC60));
  VFA U60 (.in_A(in_A[60]), .in_B(in_B[60]), .in_CI(nC60), .out_S(out_S[60]), .out_CO(nC61));
  VFA U61 (.in_A(in_A[61]), .in_B(in_B[61]), .in_CI(nC61), .out_S(out_S[61]), .out_CO(nC62));
  VFA U62 (.in_A(in_A[62]), .in_B(in_B[62]), .in_CI(nC62), .out_S(out_S[62]), .out_CO(nC63));
  VFA U63 (.in_A(in_A[63]), .in_B(in_B[63]), .in_CI(nC63), .out_S(out_S[63]), .out_CO(nC64));
  VFA U64 (.in_A(in_A[64]), .in_B(in_B[64]), .in_CI(nC64), .out_S(out_S[64]), .out_CO(nC65));
  VFA U65 (.in_A(in_A[65]), .in_B(in_B[65]), .in_CI(nC65), .out_S(out_S[65]), .out_CO(nC66));
  VFA U66 (.in_A(in_A[66]), .in_B(in_B[66]), .in_CI(nC66), .out_S(out_S[66]), .out_CO(nC67));
  VFA U67 (.in_A(in_A[67]), .in_B(in_B[67]), .in_CI(nC67), .out_S(out_S[67]), .out_CO(nC68));
  VFA U68 (.in_A(in_A[68]), .in_B(in_B[68]), .in_CI(nC68), .out_S(out_S[68]), .out_CO(nC69));
  VFA U69 (.in_A(in_A[69]), .in_B(in_B[69]), .in_CI(nC69), .out_S(out_S[69]), .out_CO(nC70));
  VFA U70 (.in_A(in_A[70]), .in_B(in_B[70]), .in_CI(nC70), .out_S(out_S[70]), .out_CO(nC71));
  VFA U71 (.in_A(in_A[71]), .in_B(in_B[71]), .in_CI(nC71), .out_S(out_S[71]), .out_CO(nC72));
  VFA U72 (.in_A(in_A[72]), .in_B(in_B[72]), .in_CI(nC72), .out_S(out_S[72]), .out_CO(nC73));
  VFA U73 (.in_A(in_A[73]), .in_B(in_B[73]), .in_CI(nC73), .out_S(out_S[73]), .out_CO(nC74));
  VFA U74 (.in_A(in_A[74]), .in_B(in_B[74]), .in_CI(nC74), .out_S(out_S[74]), .out_CO(nC75));
  VFA U75 (.in_A(in_A[75]), .in_B(in_B[75]), .in_CI(nC75), .out_S(out_S[75]), .out_CO(nC76));
  VFA U76 (.in_A(in_A[76]), .in_B(in_B[76]), .in_CI(nC76), .out_S(out_S[76]), .out_CO(nC77));
  VFA U77 (.in_A(in_A[77]), .in_B(in_B[77]), .in_CI(nC77), .out_S(out_S[77]), .out_CO(nC78));
  VFA U78 (.in_A(in_A[78]), .in_B(in_B[78]), .in_CI(nC78), .out_S(out_S[78]), .out_CO(nC79));
  VFA U79 (.in_A(in_A[79]), .in_B(in_B[79]), .in_CI(nC79), .out_S(out_S[79]), .out_CO(nC80));
  VFA U80 (.in_A(in_A[80]), .in_B(in_B[80]), .in_CI(nC80), .out_S(out_S[80]), .out_CO(nC81));
  VFA U81 (.in_A(in_A[81]), .in_B(in_B[81]), .in_CI(nC81), .out_S(out_S[81]), .out_CO(nC82));
  VFA U82 (.in_A(in_A[82]), .in_B(in_B[82]), .in_CI(nC82), .out_S(out_S[82]), .out_CO(nC83));
  VFA U83 (.in_A(in_A[83]), .in_B(in_B[83]), .in_CI(nC83), .out_S(out_S[83]), .out_CO(nC84));
  VFA U84 (.in_A(in_A[84]), .in_B(in_B[84]), .in_CI(nC84), .out_S(out_S[84]), .out_CO(nC85));
  VFA U85 (.in_A(in_A[85]), .in_B(in_B[85]), .in_CI(nC85), .out_S(out_S[85]), .out_CO(nC86));
  VFA U86 (.in_A(in_A[86]), .in_B(in_B[86]), .in_CI(nC86), .out_S(out_S[86]), .out_CO(nC87));
  VFA U87 (.in_A(in_A[87]), .in_B(in_B[87]), .in_CI(nC87), .out_S(out_S[87]), .out_CO(nC88));
  VFA U88 (.in_A(in_A[88]), .in_B(in_B[88]), .in_CI(nC88), .out_S(out_S[88]), .out_CO(nC89));
  VFA U89 (.in_A(in_A[89]), .in_B(in_B[89]), .in_CI(nC89), .out_S(out_S[89]), .out_CO(nC90));
  VFA U90 (.in_A(in_A[90]), .in_B(in_B[90]), .in_CI(nC90), .out_S(out_S[90]), .out_CO(nC91));
  VFA U91 (.in_A(in_A[91]), .in_B(in_B[91]), .in_CI(nC91), .out_S(out_S[91]), .out_CO(nC92));
  VFA U92 (.in_A(in_A[92]), .in_B(in_B[92]), .in_CI(nC92), .out_S(out_S[92]), .out_CO(nC93));
  VFA U93 (.in_A(in_A[93]), .in_B(in_B[93]), .in_CI(nC93), .out_S(out_S[93]), .out_CO(nC94));
  VFA U94 (.in_A(in_A[94]), .in_B(in_B[94]), .in_CI(nC94), .out_S(out_S[94]), .out_CO(nC95));
  VFA U95 (.in_A(in_A[95]), .in_B(in_B[95]), .in_CI(nC95), .out_S(out_S[95]), .out_CO(nC96));
  VFA U96 (.in_A(in_A[96]), .in_B(in_B[96]), .in_CI(nC96), .out_S(out_S[96]), .out_CO(nC97));
  VFA U97 (.in_A(in_A[97]), .in_B(in_B[97]), .in_CI(nC97), .out_S(out_S[97]), .out_CO(nC98));
  VFA U98 (.in_A(in_A[98]), .in_B(in_B[98]), .in_CI(nC98), .out_S(out_S[98]), .out_CO(nC99));
  VFA U99 (.in_A(in_A[99]), .in_B(in_B[99]), .in_CI(nC99), .out_S(out_S[99]), .out_CO(nC100));
  VFA U100 (.in_A(in_A[100]), .in_B(in_B[100]), .in_CI(nC100), .out_S(out_S[100]), .out_CO(nC101));
  VFA U101 (.in_A(in_A[101]), .in_B(in_B[101]), .in_CI(nC101), .out_S(out_S[101]), .out_CO(nC102));
  VFA U102 (.in_A(in_A[102]), .in_B(in_B[102]), .in_CI(nC102), .out_S(out_S[102]), .out_CO(nC103));
  VFA U103 (.in_A(in_A[103]), .in_B(in_B[103]), .in_CI(nC103), .out_S(out_S[103]), .out_CO(nC104));
  VFA U104 (.in_A(in_A[104]), .in_B(in_B[104]), .in_CI(nC104), .out_S(out_S[104]), .out_CO(nC105));
  VFA U105 (.in_A(in_A[105]), .in_B(in_B[105]), .in_CI(nC105), .out_S(out_S[105]), .out_CO(nC106));
  VFA U106 (.in_A(in_A[106]), .in_B(in_B[106]), .in_CI(nC106), .out_S(out_S[106]), .out_CO(nC107));
  VFA U107 (.in_A(in_A[107]), .in_B(in_B[107]), .in_CI(nC107), .out_S(out_S[107]), .out_CO(nC108));
  VFA U108 (.in_A(in_A[108]), .in_B(in_B[108]), .in_CI(nC108), .out_S(out_S[108]), .out_CO(nC109));
  VFA U109 (.in_A(in_A[109]), .in_B(in_B[109]), .in_CI(nC109), .out_S(out_S[109]), .out_CO(nC110));
  VFA U110 (.in_A(in_A[110]), .in_B(in_B[110]), .in_CI(nC110), .out_S(out_S[110]), .out_CO(nC111));
  VFA U111 (.in_A(in_A[111]), .in_B(in_B[111]), .in_CI(nC111), .out_S(out_S[111]), .out_CO(nC112));
  VFA U112 (.in_A(in_A[112]), .in_B(in_B[112]), .in_CI(nC112), .out_S(out_S[112]), .out_CO(nC113));
  VFA U113 (.in_A(in_A[113]), .in_B(in_B[113]), .in_CI(nC113), .out_S(out_S[113]), .out_CO(nC114));
  VFA U114 (.in_A(in_A[114]), .in_B(in_B[114]), .in_CI(nC114), .out_S(out_S[114]), .out_CO(nC115));
  VFA U115 (.in_A(in_A[115]), .in_B(in_B[115]), .in_CI(nC115), .out_S(out_S[115]), .out_CO(nC116));
  VFA U116 (.in_A(in_A[116]), .in_B(in_B[116]), .in_CI(nC116), .out_S(out_S[116]), .out_CO(nC117));
  VFA U117 (.in_A(in_A[117]), .in_B(in_B[117]), .in_CI(nC117), .out_S(out_S[117]), .out_CO(nC118));
  VFA U118 (.in_A(in_A[118]), .in_B(in_B[118]), .in_CI(nC118), .out_S(out_S[118]), .out_CO(nC119));
  VFA U119 (.in_A(in_A[119]), .in_B(in_B[119]), .in_CI(nC119), .out_S(out_S[119]), .out_CO(nC120));
  VFA U120 (.in_A(in_A[120]), .in_B(in_B[120]), .in_CI(nC120), .out_S(out_S[120]), .out_CO(nC121));
  VFA U121 (.in_A(in_A[121]), .in_B(in_B[121]), .in_CI(nC121), .out_S(out_S[121]), .out_CO(nC122));
  VFA U122 (.in_A(in_A[122]), .in_B(in_B[122]), .in_CI(nC122), .out_S(out_S[122]), .out_CO(nC123));
  VFA U123 (.in_A(in_A[123]), .in_B(in_B[123]), .in_CI(nC123), .out_S(out_S[123]), .out_CO(nC124));
  VFA U124 (.in_A(in_A[124]), .in_B(in_B[124]), .in_CI(nC124), .out_S(out_S[124]), .out_CO(nC125));
  VFA U125 (.in_A(in_A[125]), .in_B(in_B[125]), .in_CI(nC125), .out_S(out_S[125]), .out_CO(nC126));
  VFA U126 (.in_A(in_A[126]), .in_B(in_B[126]), .in_CI(nC126), .out_S(out_S[126]), .out_CO(nC127));
  VFA U127 (.in_A(in_A[127]), .in_B(in_B[127]), .in_CI(nC127), .out_S(out_S[127]), .out_CO(out_CO));
endmodule

