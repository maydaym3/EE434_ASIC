/net/ugrads/jtschir1/pvt/ee434/tut_Innovus/lib/lef/NangateOpenCellLibrary.lef