module VHA (in_A, in_B, out_S, out_CO);
  input in_A, in_B;
  output out_S, out_CO;

  assign out_S = in_A ^ in_B;
  assign out_CO = in_A & in_B;
endmodule

module VFA (in_A, in_B, in_CI, out_S, out_CO);
  input in_A, in_B, in_CI;
  output out_S, out_CO;

  assign out_S = in_A ^ in_B ^ in_CI;
  assign out_CO = (in_A & in_B) | (in_B & in_CI) | (in_CI & in_A);
endmodule



module VCondSumAdder_64 (in_A, in_B, in_CI, out_S, out_CO);
  input [63:0] in_A, in_B;
  input in_CI;
  output [63:0] out_S;
  output out_CO;

  VHA U_st1_b0_c0 (.in_A(in_A[0]), .in_B(in_B[0]), .out_S(nS_st1_b0_c0), .out_CO(nC_st1_b0_c0));
  VFA U_st1_b0_c1 (.in_A(in_A[0]), .in_B(in_B[0]), .in_CI(1'b1), .out_S(nS_st1_b0_c1), .out_CO(nC_st1_b0_c1));
  VHA U_st1_b1_c0 (.in_A(in_A[1]), .in_B(in_B[1]), .out_S(nS_st1_b1_c0), .out_CO(nC_st1_b1_c0));
  VFA U_st1_b1_c1 (.in_A(in_A[1]), .in_B(in_B[1]), .in_CI(1'b1), .out_S(nS_st1_b1_c1), .out_CO(nC_st1_b1_c1));
  VHA U_st1_b2_c0 (.in_A(in_A[2]), .in_B(in_B[2]), .out_S(nS_st1_b2_c0), .out_CO(nC_st1_b2_c0));
  VFA U_st1_b2_c1 (.in_A(in_A[2]), .in_B(in_B[2]), .in_CI(1'b1), .out_S(nS_st1_b2_c1), .out_CO(nC_st1_b2_c1));
  VHA U_st1_b3_c0 (.in_A(in_A[3]), .in_B(in_B[3]), .out_S(nS_st1_b3_c0), .out_CO(nC_st1_b3_c0));
  VFA U_st1_b3_c1 (.in_A(in_A[3]), .in_B(in_B[3]), .in_CI(1'b1), .out_S(nS_st1_b3_c1), .out_CO(nC_st1_b3_c1));
  VHA U_st1_b4_c0 (.in_A(in_A[4]), .in_B(in_B[4]), .out_S(nS_st1_b4_c0), .out_CO(nC_st1_b4_c0));
  VFA U_st1_b4_c1 (.in_A(in_A[4]), .in_B(in_B[4]), .in_CI(1'b1), .out_S(nS_st1_b4_c1), .out_CO(nC_st1_b4_c1));
  VHA U_st1_b5_c0 (.in_A(in_A[5]), .in_B(in_B[5]), .out_S(nS_st1_b5_c0), .out_CO(nC_st1_b5_c0));
  VFA U_st1_b5_c1 (.in_A(in_A[5]), .in_B(in_B[5]), .in_CI(1'b1), .out_S(nS_st1_b5_c1), .out_CO(nC_st1_b5_c1));
  VHA U_st1_b6_c0 (.in_A(in_A[6]), .in_B(in_B[6]), .out_S(nS_st1_b6_c0), .out_CO(nC_st1_b6_c0));
  VFA U_st1_b6_c1 (.in_A(in_A[6]), .in_B(in_B[6]), .in_CI(1'b1), .out_S(nS_st1_b6_c1), .out_CO(nC_st1_b6_c1));
  VHA U_st1_b7_c0 (.in_A(in_A[7]), .in_B(in_B[7]), .out_S(nS_st1_b7_c0), .out_CO(nC_st1_b7_c0));
  VFA U_st1_b7_c1 (.in_A(in_A[7]), .in_B(in_B[7]), .in_CI(1'b1), .out_S(nS_st1_b7_c1), .out_CO(nC_st1_b7_c1));
  VHA U_st1_b8_c0 (.in_A(in_A[8]), .in_B(in_B[8]), .out_S(nS_st1_b8_c0), .out_CO(nC_st1_b8_c0));
  VFA U_st1_b8_c1 (.in_A(in_A[8]), .in_B(in_B[8]), .in_CI(1'b1), .out_S(nS_st1_b8_c1), .out_CO(nC_st1_b8_c1));
  VHA U_st1_b9_c0 (.in_A(in_A[9]), .in_B(in_B[9]), .out_S(nS_st1_b9_c0), .out_CO(nC_st1_b9_c0));
  VFA U_st1_b9_c1 (.in_A(in_A[9]), .in_B(in_B[9]), .in_CI(1'b1), .out_S(nS_st1_b9_c1), .out_CO(nC_st1_b9_c1));
  VHA U_st1_b10_c0 (.in_A(in_A[10]), .in_B(in_B[10]), .out_S(nS_st1_b10_c0), .out_CO(nC_st1_b10_c0));
  VFA U_st1_b10_c1 (.in_A(in_A[10]), .in_B(in_B[10]), .in_CI(1'b1), .out_S(nS_st1_b10_c1), .out_CO(nC_st1_b10_c1));
  VHA U_st1_b11_c0 (.in_A(in_A[11]), .in_B(in_B[11]), .out_S(nS_st1_b11_c0), .out_CO(nC_st1_b11_c0));
  VFA U_st1_b11_c1 (.in_A(in_A[11]), .in_B(in_B[11]), .in_CI(1'b1), .out_S(nS_st1_b11_c1), .out_CO(nC_st1_b11_c1));
  VHA U_st1_b12_c0 (.in_A(in_A[12]), .in_B(in_B[12]), .out_S(nS_st1_b12_c0), .out_CO(nC_st1_b12_c0));
  VFA U_st1_b12_c1 (.in_A(in_A[12]), .in_B(in_B[12]), .in_CI(1'b1), .out_S(nS_st1_b12_c1), .out_CO(nC_st1_b12_c1));
  VHA U_st1_b13_c0 (.in_A(in_A[13]), .in_B(in_B[13]), .out_S(nS_st1_b13_c0), .out_CO(nC_st1_b13_c0));
  VFA U_st1_b13_c1 (.in_A(in_A[13]), .in_B(in_B[13]), .in_CI(1'b1), .out_S(nS_st1_b13_c1), .out_CO(nC_st1_b13_c1));
  VHA U_st1_b14_c0 (.in_A(in_A[14]), .in_B(in_B[14]), .out_S(nS_st1_b14_c0), .out_CO(nC_st1_b14_c0));
  VFA U_st1_b14_c1 (.in_A(in_A[14]), .in_B(in_B[14]), .in_CI(1'b1), .out_S(nS_st1_b14_c1), .out_CO(nC_st1_b14_c1));
  VHA U_st1_b15_c0 (.in_A(in_A[15]), .in_B(in_B[15]), .out_S(nS_st1_b15_c0), .out_CO(nC_st1_b15_c0));
  VFA U_st1_b15_c1 (.in_A(in_A[15]), .in_B(in_B[15]), .in_CI(1'b1), .out_S(nS_st1_b15_c1), .out_CO(nC_st1_b15_c1));
  VHA U_st1_b16_c0 (.in_A(in_A[16]), .in_B(in_B[16]), .out_S(nS_st1_b16_c0), .out_CO(nC_st1_b16_c0));
  VFA U_st1_b16_c1 (.in_A(in_A[16]), .in_B(in_B[16]), .in_CI(1'b1), .out_S(nS_st1_b16_c1), .out_CO(nC_st1_b16_c1));
  VHA U_st1_b17_c0 (.in_A(in_A[17]), .in_B(in_B[17]), .out_S(nS_st1_b17_c0), .out_CO(nC_st1_b17_c0));
  VFA U_st1_b17_c1 (.in_A(in_A[17]), .in_B(in_B[17]), .in_CI(1'b1), .out_S(nS_st1_b17_c1), .out_CO(nC_st1_b17_c1));
  VHA U_st1_b18_c0 (.in_A(in_A[18]), .in_B(in_B[18]), .out_S(nS_st1_b18_c0), .out_CO(nC_st1_b18_c0));
  VFA U_st1_b18_c1 (.in_A(in_A[18]), .in_B(in_B[18]), .in_CI(1'b1), .out_S(nS_st1_b18_c1), .out_CO(nC_st1_b18_c1));
  VHA U_st1_b19_c0 (.in_A(in_A[19]), .in_B(in_B[19]), .out_S(nS_st1_b19_c0), .out_CO(nC_st1_b19_c0));
  VFA U_st1_b19_c1 (.in_A(in_A[19]), .in_B(in_B[19]), .in_CI(1'b1), .out_S(nS_st1_b19_c1), .out_CO(nC_st1_b19_c1));
  VHA U_st1_b20_c0 (.in_A(in_A[20]), .in_B(in_B[20]), .out_S(nS_st1_b20_c0), .out_CO(nC_st1_b20_c0));
  VFA U_st1_b20_c1 (.in_A(in_A[20]), .in_B(in_B[20]), .in_CI(1'b1), .out_S(nS_st1_b20_c1), .out_CO(nC_st1_b20_c1));
  VHA U_st1_b21_c0 (.in_A(in_A[21]), .in_B(in_B[21]), .out_S(nS_st1_b21_c0), .out_CO(nC_st1_b21_c0));
  VFA U_st1_b21_c1 (.in_A(in_A[21]), .in_B(in_B[21]), .in_CI(1'b1), .out_S(nS_st1_b21_c1), .out_CO(nC_st1_b21_c1));
  VHA U_st1_b22_c0 (.in_A(in_A[22]), .in_B(in_B[22]), .out_S(nS_st1_b22_c0), .out_CO(nC_st1_b22_c0));
  VFA U_st1_b22_c1 (.in_A(in_A[22]), .in_B(in_B[22]), .in_CI(1'b1), .out_S(nS_st1_b22_c1), .out_CO(nC_st1_b22_c1));
  VHA U_st1_b23_c0 (.in_A(in_A[23]), .in_B(in_B[23]), .out_S(nS_st1_b23_c0), .out_CO(nC_st1_b23_c0));
  VFA U_st1_b23_c1 (.in_A(in_A[23]), .in_B(in_B[23]), .in_CI(1'b1), .out_S(nS_st1_b23_c1), .out_CO(nC_st1_b23_c1));
  VHA U_st1_b24_c0 (.in_A(in_A[24]), .in_B(in_B[24]), .out_S(nS_st1_b24_c0), .out_CO(nC_st1_b24_c0));
  VFA U_st1_b24_c1 (.in_A(in_A[24]), .in_B(in_B[24]), .in_CI(1'b1), .out_S(nS_st1_b24_c1), .out_CO(nC_st1_b24_c1));
  VHA U_st1_b25_c0 (.in_A(in_A[25]), .in_B(in_B[25]), .out_S(nS_st1_b25_c0), .out_CO(nC_st1_b25_c0));
  VFA U_st1_b25_c1 (.in_A(in_A[25]), .in_B(in_B[25]), .in_CI(1'b1), .out_S(nS_st1_b25_c1), .out_CO(nC_st1_b25_c1));
  VHA U_st1_b26_c0 (.in_A(in_A[26]), .in_B(in_B[26]), .out_S(nS_st1_b26_c0), .out_CO(nC_st1_b26_c0));
  VFA U_st1_b26_c1 (.in_A(in_A[26]), .in_B(in_B[26]), .in_CI(1'b1), .out_S(nS_st1_b26_c1), .out_CO(nC_st1_b26_c1));
  VHA U_st1_b27_c0 (.in_A(in_A[27]), .in_B(in_B[27]), .out_S(nS_st1_b27_c0), .out_CO(nC_st1_b27_c0));
  VFA U_st1_b27_c1 (.in_A(in_A[27]), .in_B(in_B[27]), .in_CI(1'b1), .out_S(nS_st1_b27_c1), .out_CO(nC_st1_b27_c1));
  VHA U_st1_b28_c0 (.in_A(in_A[28]), .in_B(in_B[28]), .out_S(nS_st1_b28_c0), .out_CO(nC_st1_b28_c0));
  VFA U_st1_b28_c1 (.in_A(in_A[28]), .in_B(in_B[28]), .in_CI(1'b1), .out_S(nS_st1_b28_c1), .out_CO(nC_st1_b28_c1));
  VHA U_st1_b29_c0 (.in_A(in_A[29]), .in_B(in_B[29]), .out_S(nS_st1_b29_c0), .out_CO(nC_st1_b29_c0));
  VFA U_st1_b29_c1 (.in_A(in_A[29]), .in_B(in_B[29]), .in_CI(1'b1), .out_S(nS_st1_b29_c1), .out_CO(nC_st1_b29_c1));
  VHA U_st1_b30_c0 (.in_A(in_A[30]), .in_B(in_B[30]), .out_S(nS_st1_b30_c0), .out_CO(nC_st1_b30_c0));
  VFA U_st1_b30_c1 (.in_A(in_A[30]), .in_B(in_B[30]), .in_CI(1'b1), .out_S(nS_st1_b30_c1), .out_CO(nC_st1_b30_c1));
  VHA U_st1_b31_c0 (.in_A(in_A[31]), .in_B(in_B[31]), .out_S(nS_st1_b31_c0), .out_CO(nC_st1_b31_c0));
  VFA U_st1_b31_c1 (.in_A(in_A[31]), .in_B(in_B[31]), .in_CI(1'b1), .out_S(nS_st1_b31_c1), .out_CO(nC_st1_b31_c1));
  VHA U_st1_b32_c0 (.in_A(in_A[32]), .in_B(in_B[32]), .out_S(nS_st1_b32_c0), .out_CO(nC_st1_b32_c0));
  VFA U_st1_b32_c1 (.in_A(in_A[32]), .in_B(in_B[32]), .in_CI(1'b1), .out_S(nS_st1_b32_c1), .out_CO(nC_st1_b32_c1));
  VHA U_st1_b33_c0 (.in_A(in_A[33]), .in_B(in_B[33]), .out_S(nS_st1_b33_c0), .out_CO(nC_st1_b33_c0));
  VFA U_st1_b33_c1 (.in_A(in_A[33]), .in_B(in_B[33]), .in_CI(1'b1), .out_S(nS_st1_b33_c1), .out_CO(nC_st1_b33_c1));
  VHA U_st1_b34_c0 (.in_A(in_A[34]), .in_B(in_B[34]), .out_S(nS_st1_b34_c0), .out_CO(nC_st1_b34_c0));
  VFA U_st1_b34_c1 (.in_A(in_A[34]), .in_B(in_B[34]), .in_CI(1'b1), .out_S(nS_st1_b34_c1), .out_CO(nC_st1_b34_c1));
  VHA U_st1_b35_c0 (.in_A(in_A[35]), .in_B(in_B[35]), .out_S(nS_st1_b35_c0), .out_CO(nC_st1_b35_c0));
  VFA U_st1_b35_c1 (.in_A(in_A[35]), .in_B(in_B[35]), .in_CI(1'b1), .out_S(nS_st1_b35_c1), .out_CO(nC_st1_b35_c1));
  VHA U_st1_b36_c0 (.in_A(in_A[36]), .in_B(in_B[36]), .out_S(nS_st1_b36_c0), .out_CO(nC_st1_b36_c0));
  VFA U_st1_b36_c1 (.in_A(in_A[36]), .in_B(in_B[36]), .in_CI(1'b1), .out_S(nS_st1_b36_c1), .out_CO(nC_st1_b36_c1));
  VHA U_st1_b37_c0 (.in_A(in_A[37]), .in_B(in_B[37]), .out_S(nS_st1_b37_c0), .out_CO(nC_st1_b37_c0));
  VFA U_st1_b37_c1 (.in_A(in_A[37]), .in_B(in_B[37]), .in_CI(1'b1), .out_S(nS_st1_b37_c1), .out_CO(nC_st1_b37_c1));
  VHA U_st1_b38_c0 (.in_A(in_A[38]), .in_B(in_B[38]), .out_S(nS_st1_b38_c0), .out_CO(nC_st1_b38_c0));
  VFA U_st1_b38_c1 (.in_A(in_A[38]), .in_B(in_B[38]), .in_CI(1'b1), .out_S(nS_st1_b38_c1), .out_CO(nC_st1_b38_c1));
  VHA U_st1_b39_c0 (.in_A(in_A[39]), .in_B(in_B[39]), .out_S(nS_st1_b39_c0), .out_CO(nC_st1_b39_c0));
  VFA U_st1_b39_c1 (.in_A(in_A[39]), .in_B(in_B[39]), .in_CI(1'b1), .out_S(nS_st1_b39_c1), .out_CO(nC_st1_b39_c1));
  VHA U_st1_b40_c0 (.in_A(in_A[40]), .in_B(in_B[40]), .out_S(nS_st1_b40_c0), .out_CO(nC_st1_b40_c0));
  VFA U_st1_b40_c1 (.in_A(in_A[40]), .in_B(in_B[40]), .in_CI(1'b1), .out_S(nS_st1_b40_c1), .out_CO(nC_st1_b40_c1));
  VHA U_st1_b41_c0 (.in_A(in_A[41]), .in_B(in_B[41]), .out_S(nS_st1_b41_c0), .out_CO(nC_st1_b41_c0));
  VFA U_st1_b41_c1 (.in_A(in_A[41]), .in_B(in_B[41]), .in_CI(1'b1), .out_S(nS_st1_b41_c1), .out_CO(nC_st1_b41_c1));
  VHA U_st1_b42_c0 (.in_A(in_A[42]), .in_B(in_B[42]), .out_S(nS_st1_b42_c0), .out_CO(nC_st1_b42_c0));
  VFA U_st1_b42_c1 (.in_A(in_A[42]), .in_B(in_B[42]), .in_CI(1'b1), .out_S(nS_st1_b42_c1), .out_CO(nC_st1_b42_c1));
  VHA U_st1_b43_c0 (.in_A(in_A[43]), .in_B(in_B[43]), .out_S(nS_st1_b43_c0), .out_CO(nC_st1_b43_c0));
  VFA U_st1_b43_c1 (.in_A(in_A[43]), .in_B(in_B[43]), .in_CI(1'b1), .out_S(nS_st1_b43_c1), .out_CO(nC_st1_b43_c1));
  VHA U_st1_b44_c0 (.in_A(in_A[44]), .in_B(in_B[44]), .out_S(nS_st1_b44_c0), .out_CO(nC_st1_b44_c0));
  VFA U_st1_b44_c1 (.in_A(in_A[44]), .in_B(in_B[44]), .in_CI(1'b1), .out_S(nS_st1_b44_c1), .out_CO(nC_st1_b44_c1));
  VHA U_st1_b45_c0 (.in_A(in_A[45]), .in_B(in_B[45]), .out_S(nS_st1_b45_c0), .out_CO(nC_st1_b45_c0));
  VFA U_st1_b45_c1 (.in_A(in_A[45]), .in_B(in_B[45]), .in_CI(1'b1), .out_S(nS_st1_b45_c1), .out_CO(nC_st1_b45_c1));
  VHA U_st1_b46_c0 (.in_A(in_A[46]), .in_B(in_B[46]), .out_S(nS_st1_b46_c0), .out_CO(nC_st1_b46_c0));
  VFA U_st1_b46_c1 (.in_A(in_A[46]), .in_B(in_B[46]), .in_CI(1'b1), .out_S(nS_st1_b46_c1), .out_CO(nC_st1_b46_c1));
  VHA U_st1_b47_c0 (.in_A(in_A[47]), .in_B(in_B[47]), .out_S(nS_st1_b47_c0), .out_CO(nC_st1_b47_c0));
  VFA U_st1_b47_c1 (.in_A(in_A[47]), .in_B(in_B[47]), .in_CI(1'b1), .out_S(nS_st1_b47_c1), .out_CO(nC_st1_b47_c1));
  VHA U_st1_b48_c0 (.in_A(in_A[48]), .in_B(in_B[48]), .out_S(nS_st1_b48_c0), .out_CO(nC_st1_b48_c0));
  VFA U_st1_b48_c1 (.in_A(in_A[48]), .in_B(in_B[48]), .in_CI(1'b1), .out_S(nS_st1_b48_c1), .out_CO(nC_st1_b48_c1));
  VHA U_st1_b49_c0 (.in_A(in_A[49]), .in_B(in_B[49]), .out_S(nS_st1_b49_c0), .out_CO(nC_st1_b49_c0));
  VFA U_st1_b49_c1 (.in_A(in_A[49]), .in_B(in_B[49]), .in_CI(1'b1), .out_S(nS_st1_b49_c1), .out_CO(nC_st1_b49_c1));
  VHA U_st1_b50_c0 (.in_A(in_A[50]), .in_B(in_B[50]), .out_S(nS_st1_b50_c0), .out_CO(nC_st1_b50_c0));
  VFA U_st1_b50_c1 (.in_A(in_A[50]), .in_B(in_B[50]), .in_CI(1'b1), .out_S(nS_st1_b50_c1), .out_CO(nC_st1_b50_c1));
  VHA U_st1_b51_c0 (.in_A(in_A[51]), .in_B(in_B[51]), .out_S(nS_st1_b51_c0), .out_CO(nC_st1_b51_c0));
  VFA U_st1_b51_c1 (.in_A(in_A[51]), .in_B(in_B[51]), .in_CI(1'b1), .out_S(nS_st1_b51_c1), .out_CO(nC_st1_b51_c1));
  VHA U_st1_b52_c0 (.in_A(in_A[52]), .in_B(in_B[52]), .out_S(nS_st1_b52_c0), .out_CO(nC_st1_b52_c0));
  VFA U_st1_b52_c1 (.in_A(in_A[52]), .in_B(in_B[52]), .in_CI(1'b1), .out_S(nS_st1_b52_c1), .out_CO(nC_st1_b52_c1));
  VHA U_st1_b53_c0 (.in_A(in_A[53]), .in_B(in_B[53]), .out_S(nS_st1_b53_c0), .out_CO(nC_st1_b53_c0));
  VFA U_st1_b53_c1 (.in_A(in_A[53]), .in_B(in_B[53]), .in_CI(1'b1), .out_S(nS_st1_b53_c1), .out_CO(nC_st1_b53_c1));
  VHA U_st1_b54_c0 (.in_A(in_A[54]), .in_B(in_B[54]), .out_S(nS_st1_b54_c0), .out_CO(nC_st1_b54_c0));
  VFA U_st1_b54_c1 (.in_A(in_A[54]), .in_B(in_B[54]), .in_CI(1'b1), .out_S(nS_st1_b54_c1), .out_CO(nC_st1_b54_c1));
  VHA U_st1_b55_c0 (.in_A(in_A[55]), .in_B(in_B[55]), .out_S(nS_st1_b55_c0), .out_CO(nC_st1_b55_c0));
  VFA U_st1_b55_c1 (.in_A(in_A[55]), .in_B(in_B[55]), .in_CI(1'b1), .out_S(nS_st1_b55_c1), .out_CO(nC_st1_b55_c1));
  VHA U_st1_b56_c0 (.in_A(in_A[56]), .in_B(in_B[56]), .out_S(nS_st1_b56_c0), .out_CO(nC_st1_b56_c0));
  VFA U_st1_b56_c1 (.in_A(in_A[56]), .in_B(in_B[56]), .in_CI(1'b1), .out_S(nS_st1_b56_c1), .out_CO(nC_st1_b56_c1));
  VHA U_st1_b57_c0 (.in_A(in_A[57]), .in_B(in_B[57]), .out_S(nS_st1_b57_c0), .out_CO(nC_st1_b57_c0));
  VFA U_st1_b57_c1 (.in_A(in_A[57]), .in_B(in_B[57]), .in_CI(1'b1), .out_S(nS_st1_b57_c1), .out_CO(nC_st1_b57_c1));
  VHA U_st1_b58_c0 (.in_A(in_A[58]), .in_B(in_B[58]), .out_S(nS_st1_b58_c0), .out_CO(nC_st1_b58_c0));
  VFA U_st1_b58_c1 (.in_A(in_A[58]), .in_B(in_B[58]), .in_CI(1'b1), .out_S(nS_st1_b58_c1), .out_CO(nC_st1_b58_c1));
  VHA U_st1_b59_c0 (.in_A(in_A[59]), .in_B(in_B[59]), .out_S(nS_st1_b59_c0), .out_CO(nC_st1_b59_c0));
  VFA U_st1_b59_c1 (.in_A(in_A[59]), .in_B(in_B[59]), .in_CI(1'b1), .out_S(nS_st1_b59_c1), .out_CO(nC_st1_b59_c1));
  VHA U_st1_b60_c0 (.in_A(in_A[60]), .in_B(in_B[60]), .out_S(nS_st1_b60_c0), .out_CO(nC_st1_b60_c0));
  VFA U_st1_b60_c1 (.in_A(in_A[60]), .in_B(in_B[60]), .in_CI(1'b1), .out_S(nS_st1_b60_c1), .out_CO(nC_st1_b60_c1));
  VHA U_st1_b61_c0 (.in_A(in_A[61]), .in_B(in_B[61]), .out_S(nS_st1_b61_c0), .out_CO(nC_st1_b61_c0));
  VFA U_st1_b61_c1 (.in_A(in_A[61]), .in_B(in_B[61]), .in_CI(1'b1), .out_S(nS_st1_b61_c1), .out_CO(nC_st1_b61_c1));
  VHA U_st1_b62_c0 (.in_A(in_A[62]), .in_B(in_B[62]), .out_S(nS_st1_b62_c0), .out_CO(nC_st1_b62_c0));
  VFA U_st1_b62_c1 (.in_A(in_A[62]), .in_B(in_B[62]), .in_CI(1'b1), .out_S(nS_st1_b62_c1), .out_CO(nC_st1_b62_c1));
  VHA U_st1_b63_c0 (.in_A(in_A[63]), .in_B(in_B[63]), .out_S(nS_st1_b63_c0), .out_CO(nC_st1_b63_c0));
  VFA U_st1_b63_c1 (.in_A(in_A[63]), .in_B(in_B[63]), .in_CI(1'b1), .out_S(nS_st1_b63_c1), .out_CO(nC_st1_b63_c1));

  assign nS_st2_b0_c0 = nS_st1_b0_c0;
  assign nS_st2_b1_c0 = (nC_st1_b0_c0 == 0) ? nS_st1_b1_c0 : nS_st1_b1_c1;
  assign nS_st2_b2_c0 = nS_st1_b2_c0;
  assign nS_st2_b3_c0 = (nC_st1_b2_c0 == 0) ? nS_st1_b3_c0 : nS_st1_b3_c1;
  assign nS_st2_b4_c0 = nS_st1_b4_c0;
  assign nS_st2_b5_c0 = (nC_st1_b4_c0 == 0) ? nS_st1_b5_c0 : nS_st1_b5_c1;
  assign nS_st2_b6_c0 = nS_st1_b6_c0;
  assign nS_st2_b7_c0 = (nC_st1_b6_c0 == 0) ? nS_st1_b7_c0 : nS_st1_b7_c1;
  assign nS_st2_b8_c0 = nS_st1_b8_c0;
  assign nS_st2_b9_c0 = (nC_st1_b8_c0 == 0) ? nS_st1_b9_c0 : nS_st1_b9_c1;
  assign nS_st2_b10_c0 = nS_st1_b10_c0;
  assign nS_st2_b11_c0 = (nC_st1_b10_c0 == 0) ? nS_st1_b11_c0 : nS_st1_b11_c1;
  assign nS_st2_b12_c0 = nS_st1_b12_c0;
  assign nS_st2_b13_c0 = (nC_st1_b12_c0 == 0) ? nS_st1_b13_c0 : nS_st1_b13_c1;
  assign nS_st2_b14_c0 = nS_st1_b14_c0;
  assign nS_st2_b15_c0 = (nC_st1_b14_c0 == 0) ? nS_st1_b15_c0 : nS_st1_b15_c1;
  assign nS_st2_b16_c0 = nS_st1_b16_c0;
  assign nS_st2_b17_c0 = (nC_st1_b16_c0 == 0) ? nS_st1_b17_c0 : nS_st1_b17_c1;
  assign nS_st2_b18_c0 = nS_st1_b18_c0;
  assign nS_st2_b19_c0 = (nC_st1_b18_c0 == 0) ? nS_st1_b19_c0 : nS_st1_b19_c1;
  assign nS_st2_b20_c0 = nS_st1_b20_c0;
  assign nS_st2_b21_c0 = (nC_st1_b20_c0 == 0) ? nS_st1_b21_c0 : nS_st1_b21_c1;
  assign nS_st2_b22_c0 = nS_st1_b22_c0;
  assign nS_st2_b23_c0 = (nC_st1_b22_c0 == 0) ? nS_st1_b23_c0 : nS_st1_b23_c1;
  assign nS_st2_b24_c0 = nS_st1_b24_c0;
  assign nS_st2_b25_c0 = (nC_st1_b24_c0 == 0) ? nS_st1_b25_c0 : nS_st1_b25_c1;
  assign nS_st2_b26_c0 = nS_st1_b26_c0;
  assign nS_st2_b27_c0 = (nC_st1_b26_c0 == 0) ? nS_st1_b27_c0 : nS_st1_b27_c1;
  assign nS_st2_b28_c0 = nS_st1_b28_c0;
  assign nS_st2_b29_c0 = (nC_st1_b28_c0 == 0) ? nS_st1_b29_c0 : nS_st1_b29_c1;
  assign nS_st2_b30_c0 = nS_st1_b30_c0;
  assign nS_st2_b31_c0 = (nC_st1_b30_c0 == 0) ? nS_st1_b31_c0 : nS_st1_b31_c1;
  assign nS_st2_b32_c0 = nS_st1_b32_c0;
  assign nS_st2_b33_c0 = (nC_st1_b32_c0 == 0) ? nS_st1_b33_c0 : nS_st1_b33_c1;
  assign nS_st2_b34_c0 = nS_st1_b34_c0;
  assign nS_st2_b35_c0 = (nC_st1_b34_c0 == 0) ? nS_st1_b35_c0 : nS_st1_b35_c1;
  assign nS_st2_b36_c0 = nS_st1_b36_c0;
  assign nS_st2_b37_c0 = (nC_st1_b36_c0 == 0) ? nS_st1_b37_c0 : nS_st1_b37_c1;
  assign nS_st2_b38_c0 = nS_st1_b38_c0;
  assign nS_st2_b39_c0 = (nC_st1_b38_c0 == 0) ? nS_st1_b39_c0 : nS_st1_b39_c1;
  assign nS_st2_b40_c0 = nS_st1_b40_c0;
  assign nS_st2_b41_c0 = (nC_st1_b40_c0 == 0) ? nS_st1_b41_c0 : nS_st1_b41_c1;
  assign nS_st2_b42_c0 = nS_st1_b42_c0;
  assign nS_st2_b43_c0 = (nC_st1_b42_c0 == 0) ? nS_st1_b43_c0 : nS_st1_b43_c1;
  assign nS_st2_b44_c0 = nS_st1_b44_c0;
  assign nS_st2_b45_c0 = (nC_st1_b44_c0 == 0) ? nS_st1_b45_c0 : nS_st1_b45_c1;
  assign nS_st2_b46_c0 = nS_st1_b46_c0;
  assign nS_st2_b47_c0 = (nC_st1_b46_c0 == 0) ? nS_st1_b47_c0 : nS_st1_b47_c1;
  assign nS_st2_b48_c0 = nS_st1_b48_c0;
  assign nS_st2_b49_c0 = (nC_st1_b48_c0 == 0) ? nS_st1_b49_c0 : nS_st1_b49_c1;
  assign nS_st2_b50_c0 = nS_st1_b50_c0;
  assign nS_st2_b51_c0 = (nC_st1_b50_c0 == 0) ? nS_st1_b51_c0 : nS_st1_b51_c1;
  assign nS_st2_b52_c0 = nS_st1_b52_c0;
  assign nS_st2_b53_c0 = (nC_st1_b52_c0 == 0) ? nS_st1_b53_c0 : nS_st1_b53_c1;
  assign nS_st2_b54_c0 = nS_st1_b54_c0;
  assign nS_st2_b55_c0 = (nC_st1_b54_c0 == 0) ? nS_st1_b55_c0 : nS_st1_b55_c1;
  assign nS_st2_b56_c0 = nS_st1_b56_c0;
  assign nS_st2_b57_c0 = (nC_st1_b56_c0 == 0) ? nS_st1_b57_c0 : nS_st1_b57_c1;
  assign nS_st2_b58_c0 = nS_st1_b58_c0;
  assign nS_st2_b59_c0 = (nC_st1_b58_c0 == 0) ? nS_st1_b59_c0 : nS_st1_b59_c1;
  assign nS_st2_b60_c0 = nS_st1_b60_c0;
  assign nS_st2_b61_c0 = (nC_st1_b60_c0 == 0) ? nS_st1_b61_c0 : nS_st1_b61_c1;
  assign nS_st2_b62_c0 = nS_st1_b62_c0;
  assign nS_st2_b63_c0 = (nC_st1_b62_c0 == 0) ? nS_st1_b63_c0 : nS_st1_b63_c1;
  assign nS_st2_b0_c1 = nS_st1_b0_c1;
  assign nS_st2_b1_c1 = (nC_st1_b0_c1 == 0) ? nS_st1_b1_c0 : nS_st1_b1_c1;
  assign nS_st2_b2_c1 = nS_st1_b2_c1;
  assign nS_st2_b3_c1 = (nC_st1_b2_c1 == 0) ? nS_st1_b3_c0 : nS_st1_b3_c1;
  assign nS_st2_b4_c1 = nS_st1_b4_c1;
  assign nS_st2_b5_c1 = (nC_st1_b4_c1 == 0) ? nS_st1_b5_c0 : nS_st1_b5_c1;
  assign nS_st2_b6_c1 = nS_st1_b6_c1;
  assign nS_st2_b7_c1 = (nC_st1_b6_c1 == 0) ? nS_st1_b7_c0 : nS_st1_b7_c1;
  assign nS_st2_b8_c1 = nS_st1_b8_c1;
  assign nS_st2_b9_c1 = (nC_st1_b8_c1 == 0) ? nS_st1_b9_c0 : nS_st1_b9_c1;
  assign nS_st2_b10_c1 = nS_st1_b10_c1;
  assign nS_st2_b11_c1 = (nC_st1_b10_c1 == 0) ? nS_st1_b11_c0 : nS_st1_b11_c1;
  assign nS_st2_b12_c1 = nS_st1_b12_c1;
  assign nS_st2_b13_c1 = (nC_st1_b12_c1 == 0) ? nS_st1_b13_c0 : nS_st1_b13_c1;
  assign nS_st2_b14_c1 = nS_st1_b14_c1;
  assign nS_st2_b15_c1 = (nC_st1_b14_c1 == 0) ? nS_st1_b15_c0 : nS_st1_b15_c1;
  assign nS_st2_b16_c1 = nS_st1_b16_c1;
  assign nS_st2_b17_c1 = (nC_st1_b16_c1 == 0) ? nS_st1_b17_c0 : nS_st1_b17_c1;
  assign nS_st2_b18_c1 = nS_st1_b18_c1;
  assign nS_st2_b19_c1 = (nC_st1_b18_c1 == 0) ? nS_st1_b19_c0 : nS_st1_b19_c1;
  assign nS_st2_b20_c1 = nS_st1_b20_c1;
  assign nS_st2_b21_c1 = (nC_st1_b20_c1 == 0) ? nS_st1_b21_c0 : nS_st1_b21_c1;
  assign nS_st2_b22_c1 = nS_st1_b22_c1;
  assign nS_st2_b23_c1 = (nC_st1_b22_c1 == 0) ? nS_st1_b23_c0 : nS_st1_b23_c1;
  assign nS_st2_b24_c1 = nS_st1_b24_c1;
  assign nS_st2_b25_c1 = (nC_st1_b24_c1 == 0) ? nS_st1_b25_c0 : nS_st1_b25_c1;
  assign nS_st2_b26_c1 = nS_st1_b26_c1;
  assign nS_st2_b27_c1 = (nC_st1_b26_c1 == 0) ? nS_st1_b27_c0 : nS_st1_b27_c1;
  assign nS_st2_b28_c1 = nS_st1_b28_c1;
  assign nS_st2_b29_c1 = (nC_st1_b28_c1 == 0) ? nS_st1_b29_c0 : nS_st1_b29_c1;
  assign nS_st2_b30_c1 = nS_st1_b30_c1;
  assign nS_st2_b31_c1 = (nC_st1_b30_c1 == 0) ? nS_st1_b31_c0 : nS_st1_b31_c1;
  assign nS_st2_b32_c1 = nS_st1_b32_c1;
  assign nS_st2_b33_c1 = (nC_st1_b32_c1 == 0) ? nS_st1_b33_c0 : nS_st1_b33_c1;
  assign nS_st2_b34_c1 = nS_st1_b34_c1;
  assign nS_st2_b35_c1 = (nC_st1_b34_c1 == 0) ? nS_st1_b35_c0 : nS_st1_b35_c1;
  assign nS_st2_b36_c1 = nS_st1_b36_c1;
  assign nS_st2_b37_c1 = (nC_st1_b36_c1 == 0) ? nS_st1_b37_c0 : nS_st1_b37_c1;
  assign nS_st2_b38_c1 = nS_st1_b38_c1;
  assign nS_st2_b39_c1 = (nC_st1_b38_c1 == 0) ? nS_st1_b39_c0 : nS_st1_b39_c1;
  assign nS_st2_b40_c1 = nS_st1_b40_c1;
  assign nS_st2_b41_c1 = (nC_st1_b40_c1 == 0) ? nS_st1_b41_c0 : nS_st1_b41_c1;
  assign nS_st2_b42_c1 = nS_st1_b42_c1;
  assign nS_st2_b43_c1 = (nC_st1_b42_c1 == 0) ? nS_st1_b43_c0 : nS_st1_b43_c1;
  assign nS_st2_b44_c1 = nS_st1_b44_c1;
  assign nS_st2_b45_c1 = (nC_st1_b44_c1 == 0) ? nS_st1_b45_c0 : nS_st1_b45_c1;
  assign nS_st2_b46_c1 = nS_st1_b46_c1;
  assign nS_st2_b47_c1 = (nC_st1_b46_c1 == 0) ? nS_st1_b47_c0 : nS_st1_b47_c1;
  assign nS_st2_b48_c1 = nS_st1_b48_c1;
  assign nS_st2_b49_c1 = (nC_st1_b48_c1 == 0) ? nS_st1_b49_c0 : nS_st1_b49_c1;
  assign nS_st2_b50_c1 = nS_st1_b50_c1;
  assign nS_st2_b51_c1 = (nC_st1_b50_c1 == 0) ? nS_st1_b51_c0 : nS_st1_b51_c1;
  assign nS_st2_b52_c1 = nS_st1_b52_c1;
  assign nS_st2_b53_c1 = (nC_st1_b52_c1 == 0) ? nS_st1_b53_c0 : nS_st1_b53_c1;
  assign nS_st2_b54_c1 = nS_st1_b54_c1;
  assign nS_st2_b55_c1 = (nC_st1_b54_c1 == 0) ? nS_st1_b55_c0 : nS_st1_b55_c1;
  assign nS_st2_b56_c1 = nS_st1_b56_c1;
  assign nS_st2_b57_c1 = (nC_st1_b56_c1 == 0) ? nS_st1_b57_c0 : nS_st1_b57_c1;
  assign nS_st2_b58_c1 = nS_st1_b58_c1;
  assign nS_st2_b59_c1 = (nC_st1_b58_c1 == 0) ? nS_st1_b59_c0 : nS_st1_b59_c1;
  assign nS_st2_b60_c1 = nS_st1_b60_c1;
  assign nS_st2_b61_c1 = (nC_st1_b60_c1 == 0) ? nS_st1_b61_c0 : nS_st1_b61_c1;
  assign nS_st2_b62_c1 = nS_st1_b62_c1;
  assign nS_st2_b63_c1 = (nC_st1_b62_c1 == 0) ? nS_st1_b63_c0 : nS_st1_b63_c1;
  assign nC_st2_b1_c0 = (nC_st1_b0_c0 == 0) ? nC_st1_b1_c0 : nC_st1_b1_c1;
  assign nC_st2_b3_c0 = (nC_st1_b2_c0 == 0) ? nC_st1_b3_c0 : nC_st1_b3_c1;
  assign nC_st2_b5_c0 = (nC_st1_b4_c0 == 0) ? nC_st1_b5_c0 : nC_st1_b5_c1;
  assign nC_st2_b7_c0 = (nC_st1_b6_c0 == 0) ? nC_st1_b7_c0 : nC_st1_b7_c1;
  assign nC_st2_b9_c0 = (nC_st1_b8_c0 == 0) ? nC_st1_b9_c0 : nC_st1_b9_c1;
  assign nC_st2_b11_c0 = (nC_st1_b10_c0 == 0) ? nC_st1_b11_c0 : nC_st1_b11_c1;
  assign nC_st2_b13_c0 = (nC_st1_b12_c0 == 0) ? nC_st1_b13_c0 : nC_st1_b13_c1;
  assign nC_st2_b15_c0 = (nC_st1_b14_c0 == 0) ? nC_st1_b15_c0 : nC_st1_b15_c1;
  assign nC_st2_b17_c0 = (nC_st1_b16_c0 == 0) ? nC_st1_b17_c0 : nC_st1_b17_c1;
  assign nC_st2_b19_c0 = (nC_st1_b18_c0 == 0) ? nC_st1_b19_c0 : nC_st1_b19_c1;
  assign nC_st2_b21_c0 = (nC_st1_b20_c0 == 0) ? nC_st1_b21_c0 : nC_st1_b21_c1;
  assign nC_st2_b23_c0 = (nC_st1_b22_c0 == 0) ? nC_st1_b23_c0 : nC_st1_b23_c1;
  assign nC_st2_b25_c0 = (nC_st1_b24_c0 == 0) ? nC_st1_b25_c0 : nC_st1_b25_c1;
  assign nC_st2_b27_c0 = (nC_st1_b26_c0 == 0) ? nC_st1_b27_c0 : nC_st1_b27_c1;
  assign nC_st2_b29_c0 = (nC_st1_b28_c0 == 0) ? nC_st1_b29_c0 : nC_st1_b29_c1;
  assign nC_st2_b31_c0 = (nC_st1_b30_c0 == 0) ? nC_st1_b31_c0 : nC_st1_b31_c1;
  assign nC_st2_b33_c0 = (nC_st1_b32_c0 == 0) ? nC_st1_b33_c0 : nC_st1_b33_c1;
  assign nC_st2_b35_c0 = (nC_st1_b34_c0 == 0) ? nC_st1_b35_c0 : nC_st1_b35_c1;
  assign nC_st2_b37_c0 = (nC_st1_b36_c0 == 0) ? nC_st1_b37_c0 : nC_st1_b37_c1;
  assign nC_st2_b39_c0 = (nC_st1_b38_c0 == 0) ? nC_st1_b39_c0 : nC_st1_b39_c1;
  assign nC_st2_b41_c0 = (nC_st1_b40_c0 == 0) ? nC_st1_b41_c0 : nC_st1_b41_c1;
  assign nC_st2_b43_c0 = (nC_st1_b42_c0 == 0) ? nC_st1_b43_c0 : nC_st1_b43_c1;
  assign nC_st2_b45_c0 = (nC_st1_b44_c0 == 0) ? nC_st1_b45_c0 : nC_st1_b45_c1;
  assign nC_st2_b47_c0 = (nC_st1_b46_c0 == 0) ? nC_st1_b47_c0 : nC_st1_b47_c1;
  assign nC_st2_b49_c0 = (nC_st1_b48_c0 == 0) ? nC_st1_b49_c0 : nC_st1_b49_c1;
  assign nC_st2_b51_c0 = (nC_st1_b50_c0 == 0) ? nC_st1_b51_c0 : nC_st1_b51_c1;
  assign nC_st2_b53_c0 = (nC_st1_b52_c0 == 0) ? nC_st1_b53_c0 : nC_st1_b53_c1;
  assign nC_st2_b55_c0 = (nC_st1_b54_c0 == 0) ? nC_st1_b55_c0 : nC_st1_b55_c1;
  assign nC_st2_b57_c0 = (nC_st1_b56_c0 == 0) ? nC_st1_b57_c0 : nC_st1_b57_c1;
  assign nC_st2_b59_c0 = (nC_st1_b58_c0 == 0) ? nC_st1_b59_c0 : nC_st1_b59_c1;
  assign nC_st2_b61_c0 = (nC_st1_b60_c0 == 0) ? nC_st1_b61_c0 : nC_st1_b61_c1;
  assign nC_st2_b63_c0 = (nC_st1_b62_c0 == 0) ? nC_st1_b63_c0 : nC_st1_b63_c1;
  assign nC_st2_b1_c1 = (nC_st1_b0_c1 == 0) ? nC_st1_b1_c0 : nC_st1_b1_c1;
  assign nC_st2_b3_c1 = (nC_st1_b2_c1 == 0) ? nC_st1_b3_c0 : nC_st1_b3_c1;
  assign nC_st2_b5_c1 = (nC_st1_b4_c1 == 0) ? nC_st1_b5_c0 : nC_st1_b5_c1;
  assign nC_st2_b7_c1 = (nC_st1_b6_c1 == 0) ? nC_st1_b7_c0 : nC_st1_b7_c1;
  assign nC_st2_b9_c1 = (nC_st1_b8_c1 == 0) ? nC_st1_b9_c0 : nC_st1_b9_c1;
  assign nC_st2_b11_c1 = (nC_st1_b10_c1 == 0) ? nC_st1_b11_c0 : nC_st1_b11_c1;
  assign nC_st2_b13_c1 = (nC_st1_b12_c1 == 0) ? nC_st1_b13_c0 : nC_st1_b13_c1;
  assign nC_st2_b15_c1 = (nC_st1_b14_c1 == 0) ? nC_st1_b15_c0 : nC_st1_b15_c1;
  assign nC_st2_b17_c1 = (nC_st1_b16_c1 == 0) ? nC_st1_b17_c0 : nC_st1_b17_c1;
  assign nC_st2_b19_c1 = (nC_st1_b18_c1 == 0) ? nC_st1_b19_c0 : nC_st1_b19_c1;
  assign nC_st2_b21_c1 = (nC_st1_b20_c1 == 0) ? nC_st1_b21_c0 : nC_st1_b21_c1;
  assign nC_st2_b23_c1 = (nC_st1_b22_c1 == 0) ? nC_st1_b23_c0 : nC_st1_b23_c1;
  assign nC_st2_b25_c1 = (nC_st1_b24_c1 == 0) ? nC_st1_b25_c0 : nC_st1_b25_c1;
  assign nC_st2_b27_c1 = (nC_st1_b26_c1 == 0) ? nC_st1_b27_c0 : nC_st1_b27_c1;
  assign nC_st2_b29_c1 = (nC_st1_b28_c1 == 0) ? nC_st1_b29_c0 : nC_st1_b29_c1;
  assign nC_st2_b31_c1 = (nC_st1_b30_c1 == 0) ? nC_st1_b31_c0 : nC_st1_b31_c1;
  assign nC_st2_b33_c1 = (nC_st1_b32_c1 == 0) ? nC_st1_b33_c0 : nC_st1_b33_c1;
  assign nC_st2_b35_c1 = (nC_st1_b34_c1 == 0) ? nC_st1_b35_c0 : nC_st1_b35_c1;
  assign nC_st2_b37_c1 = (nC_st1_b36_c1 == 0) ? nC_st1_b37_c0 : nC_st1_b37_c1;
  assign nC_st2_b39_c1 = (nC_st1_b38_c1 == 0) ? nC_st1_b39_c0 : nC_st1_b39_c1;
  assign nC_st2_b41_c1 = (nC_st1_b40_c1 == 0) ? nC_st1_b41_c0 : nC_st1_b41_c1;
  assign nC_st2_b43_c1 = (nC_st1_b42_c1 == 0) ? nC_st1_b43_c0 : nC_st1_b43_c1;
  assign nC_st2_b45_c1 = (nC_st1_b44_c1 == 0) ? nC_st1_b45_c0 : nC_st1_b45_c1;
  assign nC_st2_b47_c1 = (nC_st1_b46_c1 == 0) ? nC_st1_b47_c0 : nC_st1_b47_c1;
  assign nC_st2_b49_c1 = (nC_st1_b48_c1 == 0) ? nC_st1_b49_c0 : nC_st1_b49_c1;
  assign nC_st2_b51_c1 = (nC_st1_b50_c1 == 0) ? nC_st1_b51_c0 : nC_st1_b51_c1;
  assign nC_st2_b53_c1 = (nC_st1_b52_c1 == 0) ? nC_st1_b53_c0 : nC_st1_b53_c1;
  assign nC_st2_b55_c1 = (nC_st1_b54_c1 == 0) ? nC_st1_b55_c0 : nC_st1_b55_c1;
  assign nC_st2_b57_c1 = (nC_st1_b56_c1 == 0) ? nC_st1_b57_c0 : nC_st1_b57_c1;
  assign nC_st2_b59_c1 = (nC_st1_b58_c1 == 0) ? nC_st1_b59_c0 : nC_st1_b59_c1;
  assign nC_st2_b61_c1 = (nC_st1_b60_c1 == 0) ? nC_st1_b61_c0 : nC_st1_b61_c1;
  assign nC_st2_b63_c1 = (nC_st1_b62_c1 == 0) ? nC_st1_b63_c0 : nC_st1_b63_c1;

  assign nS_st3_b0_c0 = nS_st2_b0_c0;
  assign nS_st3_b1_c0 = nS_st2_b1_c0;
  assign nS_st3_b2_c0 = (nC_st2_b1_c0 == 0) ? nS_st2_b2_c0 : nS_st2_b2_c1;
  assign nS_st3_b3_c0 = (nC_st2_b1_c0 == 0) ? nS_st2_b3_c0 : nS_st2_b3_c1;
  assign nS_st3_b4_c0 = nS_st2_b4_c0;
  assign nS_st3_b5_c0 = nS_st2_b5_c0;
  assign nS_st3_b6_c0 = (nC_st2_b5_c0 == 0) ? nS_st2_b6_c0 : nS_st2_b6_c1;
  assign nS_st3_b7_c0 = (nC_st2_b5_c0 == 0) ? nS_st2_b7_c0 : nS_st2_b7_c1;
  assign nS_st3_b8_c0 = nS_st2_b8_c0;
  assign nS_st3_b9_c0 = nS_st2_b9_c0;
  assign nS_st3_b10_c0 = (nC_st2_b9_c0 == 0) ? nS_st2_b10_c0 : nS_st2_b10_c1;
  assign nS_st3_b11_c0 = (nC_st2_b9_c0 == 0) ? nS_st2_b11_c0 : nS_st2_b11_c1;
  assign nS_st3_b12_c0 = nS_st2_b12_c0;
  assign nS_st3_b13_c0 = nS_st2_b13_c0;
  assign nS_st3_b14_c0 = (nC_st2_b13_c0 == 0) ? nS_st2_b14_c0 : nS_st2_b14_c1;
  assign nS_st3_b15_c0 = (nC_st2_b13_c0 == 0) ? nS_st2_b15_c0 : nS_st2_b15_c1;
  assign nS_st3_b16_c0 = nS_st2_b16_c0;
  assign nS_st3_b17_c0 = nS_st2_b17_c0;
  assign nS_st3_b18_c0 = (nC_st2_b17_c0 == 0) ? nS_st2_b18_c0 : nS_st2_b18_c1;
  assign nS_st3_b19_c0 = (nC_st2_b17_c0 == 0) ? nS_st2_b19_c0 : nS_st2_b19_c1;
  assign nS_st3_b20_c0 = nS_st2_b20_c0;
  assign nS_st3_b21_c0 = nS_st2_b21_c0;
  assign nS_st3_b22_c0 = (nC_st2_b21_c0 == 0) ? nS_st2_b22_c0 : nS_st2_b22_c1;
  assign nS_st3_b23_c0 = (nC_st2_b21_c0 == 0) ? nS_st2_b23_c0 : nS_st2_b23_c1;
  assign nS_st3_b24_c0 = nS_st2_b24_c0;
  assign nS_st3_b25_c0 = nS_st2_b25_c0;
  assign nS_st3_b26_c0 = (nC_st2_b25_c0 == 0) ? nS_st2_b26_c0 : nS_st2_b26_c1;
  assign nS_st3_b27_c0 = (nC_st2_b25_c0 == 0) ? nS_st2_b27_c0 : nS_st2_b27_c1;
  assign nS_st3_b28_c0 = nS_st2_b28_c0;
  assign nS_st3_b29_c0 = nS_st2_b29_c0;
  assign nS_st3_b30_c0 = (nC_st2_b29_c0 == 0) ? nS_st2_b30_c0 : nS_st2_b30_c1;
  assign nS_st3_b31_c0 = (nC_st2_b29_c0 == 0) ? nS_st2_b31_c0 : nS_st2_b31_c1;
  assign nS_st3_b32_c0 = nS_st2_b32_c0;
  assign nS_st3_b33_c0 = nS_st2_b33_c0;
  assign nS_st3_b34_c0 = (nC_st2_b33_c0 == 0) ? nS_st2_b34_c0 : nS_st2_b34_c1;
  assign nS_st3_b35_c0 = (nC_st2_b33_c0 == 0) ? nS_st2_b35_c0 : nS_st2_b35_c1;
  assign nS_st3_b36_c0 = nS_st2_b36_c0;
  assign nS_st3_b37_c0 = nS_st2_b37_c0;
  assign nS_st3_b38_c0 = (nC_st2_b37_c0 == 0) ? nS_st2_b38_c0 : nS_st2_b38_c1;
  assign nS_st3_b39_c0 = (nC_st2_b37_c0 == 0) ? nS_st2_b39_c0 : nS_st2_b39_c1;
  assign nS_st3_b40_c0 = nS_st2_b40_c0;
  assign nS_st3_b41_c0 = nS_st2_b41_c0;
  assign nS_st3_b42_c0 = (nC_st2_b41_c0 == 0) ? nS_st2_b42_c0 : nS_st2_b42_c1;
  assign nS_st3_b43_c0 = (nC_st2_b41_c0 == 0) ? nS_st2_b43_c0 : nS_st2_b43_c1;
  assign nS_st3_b44_c0 = nS_st2_b44_c0;
  assign nS_st3_b45_c0 = nS_st2_b45_c0;
  assign nS_st3_b46_c0 = (nC_st2_b45_c0 == 0) ? nS_st2_b46_c0 : nS_st2_b46_c1;
  assign nS_st3_b47_c0 = (nC_st2_b45_c0 == 0) ? nS_st2_b47_c0 : nS_st2_b47_c1;
  assign nS_st3_b48_c0 = nS_st2_b48_c0;
  assign nS_st3_b49_c0 = nS_st2_b49_c0;
  assign nS_st3_b50_c0 = (nC_st2_b49_c0 == 0) ? nS_st2_b50_c0 : nS_st2_b50_c1;
  assign nS_st3_b51_c0 = (nC_st2_b49_c0 == 0) ? nS_st2_b51_c0 : nS_st2_b51_c1;
  assign nS_st3_b52_c0 = nS_st2_b52_c0;
  assign nS_st3_b53_c0 = nS_st2_b53_c0;
  assign nS_st3_b54_c0 = (nC_st2_b53_c0 == 0) ? nS_st2_b54_c0 : nS_st2_b54_c1;
  assign nS_st3_b55_c0 = (nC_st2_b53_c0 == 0) ? nS_st2_b55_c0 : nS_st2_b55_c1;
  assign nS_st3_b56_c0 = nS_st2_b56_c0;
  assign nS_st3_b57_c0 = nS_st2_b57_c0;
  assign nS_st3_b58_c0 = (nC_st2_b57_c0 == 0) ? nS_st2_b58_c0 : nS_st2_b58_c1;
  assign nS_st3_b59_c0 = (nC_st2_b57_c0 == 0) ? nS_st2_b59_c0 : nS_st2_b59_c1;
  assign nS_st3_b60_c0 = nS_st2_b60_c0;
  assign nS_st3_b61_c0 = nS_st2_b61_c0;
  assign nS_st3_b62_c0 = (nC_st2_b61_c0 == 0) ? nS_st2_b62_c0 : nS_st2_b62_c1;
  assign nS_st3_b63_c0 = (nC_st2_b61_c0 == 0) ? nS_st2_b63_c0 : nS_st2_b63_c1;
  assign nS_st3_b0_c1 = nS_st2_b0_c1;
  assign nS_st3_b1_c1 = nS_st2_b1_c1;
  assign nS_st3_b2_c1 = (nC_st2_b1_c1 == 0) ? nS_st2_b2_c0 : nS_st2_b2_c1;
  assign nS_st3_b3_c1 = (nC_st2_b1_c1 == 0) ? nS_st2_b3_c0 : nS_st2_b3_c1;
  assign nS_st3_b4_c1 = nS_st2_b4_c1;
  assign nS_st3_b5_c1 = nS_st2_b5_c1;
  assign nS_st3_b6_c1 = (nC_st2_b5_c1 == 0) ? nS_st2_b6_c0 : nS_st2_b6_c1;
  assign nS_st3_b7_c1 = (nC_st2_b5_c1 == 0) ? nS_st2_b7_c0 : nS_st2_b7_c1;
  assign nS_st3_b8_c1 = nS_st2_b8_c1;
  assign nS_st3_b9_c1 = nS_st2_b9_c1;
  assign nS_st3_b10_c1 = (nC_st2_b9_c1 == 0) ? nS_st2_b10_c0 : nS_st2_b10_c1;
  assign nS_st3_b11_c1 = (nC_st2_b9_c1 == 0) ? nS_st2_b11_c0 : nS_st2_b11_c1;
  assign nS_st3_b12_c1 = nS_st2_b12_c1;
  assign nS_st3_b13_c1 = nS_st2_b13_c1;
  assign nS_st3_b14_c1 = (nC_st2_b13_c1 == 0) ? nS_st2_b14_c0 : nS_st2_b14_c1;
  assign nS_st3_b15_c1 = (nC_st2_b13_c1 == 0) ? nS_st2_b15_c0 : nS_st2_b15_c1;
  assign nS_st3_b16_c1 = nS_st2_b16_c1;
  assign nS_st3_b17_c1 = nS_st2_b17_c1;
  assign nS_st3_b18_c1 = (nC_st2_b17_c1 == 0) ? nS_st2_b18_c0 : nS_st2_b18_c1;
  assign nS_st3_b19_c1 = (nC_st2_b17_c1 == 0) ? nS_st2_b19_c0 : nS_st2_b19_c1;
  assign nS_st3_b20_c1 = nS_st2_b20_c1;
  assign nS_st3_b21_c1 = nS_st2_b21_c1;
  assign nS_st3_b22_c1 = (nC_st2_b21_c1 == 0) ? nS_st2_b22_c0 : nS_st2_b22_c1;
  assign nS_st3_b23_c1 = (nC_st2_b21_c1 == 0) ? nS_st2_b23_c0 : nS_st2_b23_c1;
  assign nS_st3_b24_c1 = nS_st2_b24_c1;
  assign nS_st3_b25_c1 = nS_st2_b25_c1;
  assign nS_st3_b26_c1 = (nC_st2_b25_c1 == 0) ? nS_st2_b26_c0 : nS_st2_b26_c1;
  assign nS_st3_b27_c1 = (nC_st2_b25_c1 == 0) ? nS_st2_b27_c0 : nS_st2_b27_c1;
  assign nS_st3_b28_c1 = nS_st2_b28_c1;
  assign nS_st3_b29_c1 = nS_st2_b29_c1;
  assign nS_st3_b30_c1 = (nC_st2_b29_c1 == 0) ? nS_st2_b30_c0 : nS_st2_b30_c1;
  assign nS_st3_b31_c1 = (nC_st2_b29_c1 == 0) ? nS_st2_b31_c0 : nS_st2_b31_c1;
  assign nS_st3_b32_c1 = nS_st2_b32_c1;
  assign nS_st3_b33_c1 = nS_st2_b33_c1;
  assign nS_st3_b34_c1 = (nC_st2_b33_c1 == 0) ? nS_st2_b34_c0 : nS_st2_b34_c1;
  assign nS_st3_b35_c1 = (nC_st2_b33_c1 == 0) ? nS_st2_b35_c0 : nS_st2_b35_c1;
  assign nS_st3_b36_c1 = nS_st2_b36_c1;
  assign nS_st3_b37_c1 = nS_st2_b37_c1;
  assign nS_st3_b38_c1 = (nC_st2_b37_c1 == 0) ? nS_st2_b38_c0 : nS_st2_b38_c1;
  assign nS_st3_b39_c1 = (nC_st2_b37_c1 == 0) ? nS_st2_b39_c0 : nS_st2_b39_c1;
  assign nS_st3_b40_c1 = nS_st2_b40_c1;
  assign nS_st3_b41_c1 = nS_st2_b41_c1;
  assign nS_st3_b42_c1 = (nC_st2_b41_c1 == 0) ? nS_st2_b42_c0 : nS_st2_b42_c1;
  assign nS_st3_b43_c1 = (nC_st2_b41_c1 == 0) ? nS_st2_b43_c0 : nS_st2_b43_c1;
  assign nS_st3_b44_c1 = nS_st2_b44_c1;
  assign nS_st3_b45_c1 = nS_st2_b45_c1;
  assign nS_st3_b46_c1 = (nC_st2_b45_c1 == 0) ? nS_st2_b46_c0 : nS_st2_b46_c1;
  assign nS_st3_b47_c1 = (nC_st2_b45_c1 == 0) ? nS_st2_b47_c0 : nS_st2_b47_c1;
  assign nS_st3_b48_c1 = nS_st2_b48_c1;
  assign nS_st3_b49_c1 = nS_st2_b49_c1;
  assign nS_st3_b50_c1 = (nC_st2_b49_c1 == 0) ? nS_st2_b50_c0 : nS_st2_b50_c1;
  assign nS_st3_b51_c1 = (nC_st2_b49_c1 == 0) ? nS_st2_b51_c0 : nS_st2_b51_c1;
  assign nS_st3_b52_c1 = nS_st2_b52_c1;
  assign nS_st3_b53_c1 = nS_st2_b53_c1;
  assign nS_st3_b54_c1 = (nC_st2_b53_c1 == 0) ? nS_st2_b54_c0 : nS_st2_b54_c1;
  assign nS_st3_b55_c1 = (nC_st2_b53_c1 == 0) ? nS_st2_b55_c0 : nS_st2_b55_c1;
  assign nS_st3_b56_c1 = nS_st2_b56_c1;
  assign nS_st3_b57_c1 = nS_st2_b57_c1;
  assign nS_st3_b58_c1 = (nC_st2_b57_c1 == 0) ? nS_st2_b58_c0 : nS_st2_b58_c1;
  assign nS_st3_b59_c1 = (nC_st2_b57_c1 == 0) ? nS_st2_b59_c0 : nS_st2_b59_c1;
  assign nS_st3_b60_c1 = nS_st2_b60_c1;
  assign nS_st3_b61_c1 = nS_st2_b61_c1;
  assign nS_st3_b62_c1 = (nC_st2_b61_c1 == 0) ? nS_st2_b62_c0 : nS_st2_b62_c1;
  assign nS_st3_b63_c1 = (nC_st2_b61_c1 == 0) ? nS_st2_b63_c0 : nS_st2_b63_c1;
  assign nC_st3_b3_c0 = (nC_st2_b1_c0 == 0) ? nC_st2_b3_c0 : nC_st2_b3_c1;
  assign nC_st3_b7_c0 = (nC_st2_b5_c0 == 0) ? nC_st2_b7_c0 : nC_st2_b7_c1;
  assign nC_st3_b11_c0 = (nC_st2_b9_c0 == 0) ? nC_st2_b11_c0 : nC_st2_b11_c1;
  assign nC_st3_b15_c0 = (nC_st2_b13_c0 == 0) ? nC_st2_b15_c0 : nC_st2_b15_c1;
  assign nC_st3_b19_c0 = (nC_st2_b17_c0 == 0) ? nC_st2_b19_c0 : nC_st2_b19_c1;
  assign nC_st3_b23_c0 = (nC_st2_b21_c0 == 0) ? nC_st2_b23_c0 : nC_st2_b23_c1;
  assign nC_st3_b27_c0 = (nC_st2_b25_c0 == 0) ? nC_st2_b27_c0 : nC_st2_b27_c1;
  assign nC_st3_b31_c0 = (nC_st2_b29_c0 == 0) ? nC_st2_b31_c0 : nC_st2_b31_c1;
  assign nC_st3_b35_c0 = (nC_st2_b33_c0 == 0) ? nC_st2_b35_c0 : nC_st2_b35_c1;
  assign nC_st3_b39_c0 = (nC_st2_b37_c0 == 0) ? nC_st2_b39_c0 : nC_st2_b39_c1;
  assign nC_st3_b43_c0 = (nC_st2_b41_c0 == 0) ? nC_st2_b43_c0 : nC_st2_b43_c1;
  assign nC_st3_b47_c0 = (nC_st2_b45_c0 == 0) ? nC_st2_b47_c0 : nC_st2_b47_c1;
  assign nC_st3_b51_c0 = (nC_st2_b49_c0 == 0) ? nC_st2_b51_c0 : nC_st2_b51_c1;
  assign nC_st3_b55_c0 = (nC_st2_b53_c0 == 0) ? nC_st2_b55_c0 : nC_st2_b55_c1;
  assign nC_st3_b59_c0 = (nC_st2_b57_c0 == 0) ? nC_st2_b59_c0 : nC_st2_b59_c1;
  assign nC_st3_b63_c0 = (nC_st2_b61_c0 == 0) ? nC_st2_b63_c0 : nC_st2_b63_c1;
  assign nC_st3_b3_c1 = (nC_st2_b1_c1 == 0) ? nC_st2_b3_c0 : nC_st2_b3_c1;
  assign nC_st3_b7_c1 = (nC_st2_b5_c1 == 0) ? nC_st2_b7_c0 : nC_st2_b7_c1;
  assign nC_st3_b11_c1 = (nC_st2_b9_c1 == 0) ? nC_st2_b11_c0 : nC_st2_b11_c1;
  assign nC_st3_b15_c1 = (nC_st2_b13_c1 == 0) ? nC_st2_b15_c0 : nC_st2_b15_c1;
  assign nC_st3_b19_c1 = (nC_st2_b17_c1 == 0) ? nC_st2_b19_c0 : nC_st2_b19_c1;
  assign nC_st3_b23_c1 = (nC_st2_b21_c1 == 0) ? nC_st2_b23_c0 : nC_st2_b23_c1;
  assign nC_st3_b27_c1 = (nC_st2_b25_c1 == 0) ? nC_st2_b27_c0 : nC_st2_b27_c1;
  assign nC_st3_b31_c1 = (nC_st2_b29_c1 == 0) ? nC_st2_b31_c0 : nC_st2_b31_c1;
  assign nC_st3_b35_c1 = (nC_st2_b33_c1 == 0) ? nC_st2_b35_c0 : nC_st2_b35_c1;
  assign nC_st3_b39_c1 = (nC_st2_b37_c1 == 0) ? nC_st2_b39_c0 : nC_st2_b39_c1;
  assign nC_st3_b43_c1 = (nC_st2_b41_c1 == 0) ? nC_st2_b43_c0 : nC_st2_b43_c1;
  assign nC_st3_b47_c1 = (nC_st2_b45_c1 == 0) ? nC_st2_b47_c0 : nC_st2_b47_c1;
  assign nC_st3_b51_c1 = (nC_st2_b49_c1 == 0) ? nC_st2_b51_c0 : nC_st2_b51_c1;
  assign nC_st3_b55_c1 = (nC_st2_b53_c1 == 0) ? nC_st2_b55_c0 : nC_st2_b55_c1;
  assign nC_st3_b59_c1 = (nC_st2_b57_c1 == 0) ? nC_st2_b59_c0 : nC_st2_b59_c1;
  assign nC_st3_b63_c1 = (nC_st2_b61_c1 == 0) ? nC_st2_b63_c0 : nC_st2_b63_c1;

  assign nS_st4_b0_c0 = nS_st3_b0_c0;
  assign nS_st4_b1_c0 = nS_st3_b1_c0;
  assign nS_st4_b2_c0 = nS_st3_b2_c0;
  assign nS_st4_b3_c0 = nS_st3_b3_c0;
  assign nS_st4_b4_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b4_c0 : nS_st3_b4_c1;
  assign nS_st4_b5_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b5_c0 : nS_st3_b5_c1;
  assign nS_st4_b6_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b6_c0 : nS_st3_b6_c1;
  assign nS_st4_b7_c0 = (nC_st3_b3_c0 == 0) ? nS_st3_b7_c0 : nS_st3_b7_c1;
  assign nS_st4_b8_c0 = nS_st3_b8_c0;
  assign nS_st4_b9_c0 = nS_st3_b9_c0;
  assign nS_st4_b10_c0 = nS_st3_b10_c0;
  assign nS_st4_b11_c0 = nS_st3_b11_c0;
  assign nS_st4_b12_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b12_c0 : nS_st3_b12_c1;
  assign nS_st4_b13_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b13_c0 : nS_st3_b13_c1;
  assign nS_st4_b14_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b14_c0 : nS_st3_b14_c1;
  assign nS_st4_b15_c0 = (nC_st3_b11_c0 == 0) ? nS_st3_b15_c0 : nS_st3_b15_c1;
  assign nS_st4_b16_c0 = nS_st3_b16_c0;
  assign nS_st4_b17_c0 = nS_st3_b17_c0;
  assign nS_st4_b18_c0 = nS_st3_b18_c0;
  assign nS_st4_b19_c0 = nS_st3_b19_c0;
  assign nS_st4_b20_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b20_c0 : nS_st3_b20_c1;
  assign nS_st4_b21_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b21_c0 : nS_st3_b21_c1;
  assign nS_st4_b22_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b22_c0 : nS_st3_b22_c1;
  assign nS_st4_b23_c0 = (nC_st3_b19_c0 == 0) ? nS_st3_b23_c0 : nS_st3_b23_c1;
  assign nS_st4_b24_c0 = nS_st3_b24_c0;
  assign nS_st4_b25_c0 = nS_st3_b25_c0;
  assign nS_st4_b26_c0 = nS_st3_b26_c0;
  assign nS_st4_b27_c0 = nS_st3_b27_c0;
  assign nS_st4_b28_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b28_c0 : nS_st3_b28_c1;
  assign nS_st4_b29_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b29_c0 : nS_st3_b29_c1;
  assign nS_st4_b30_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b30_c0 : nS_st3_b30_c1;
  assign nS_st4_b31_c0 = (nC_st3_b27_c0 == 0) ? nS_st3_b31_c0 : nS_st3_b31_c1;
  assign nS_st4_b32_c0 = nS_st3_b32_c0;
  assign nS_st4_b33_c0 = nS_st3_b33_c0;
  assign nS_st4_b34_c0 = nS_st3_b34_c0;
  assign nS_st4_b35_c0 = nS_st3_b35_c0;
  assign nS_st4_b36_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b36_c0 : nS_st3_b36_c1;
  assign nS_st4_b37_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b37_c0 : nS_st3_b37_c1;
  assign nS_st4_b38_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b38_c0 : nS_st3_b38_c1;
  assign nS_st4_b39_c0 = (nC_st3_b35_c0 == 0) ? nS_st3_b39_c0 : nS_st3_b39_c1;
  assign nS_st4_b40_c0 = nS_st3_b40_c0;
  assign nS_st4_b41_c0 = nS_st3_b41_c0;
  assign nS_st4_b42_c0 = nS_st3_b42_c0;
  assign nS_st4_b43_c0 = nS_st3_b43_c0;
  assign nS_st4_b44_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b44_c0 : nS_st3_b44_c1;
  assign nS_st4_b45_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b45_c0 : nS_st3_b45_c1;
  assign nS_st4_b46_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b46_c0 : nS_st3_b46_c1;
  assign nS_st4_b47_c0 = (nC_st3_b43_c0 == 0) ? nS_st3_b47_c0 : nS_st3_b47_c1;
  assign nS_st4_b48_c0 = nS_st3_b48_c0;
  assign nS_st4_b49_c0 = nS_st3_b49_c0;
  assign nS_st4_b50_c0 = nS_st3_b50_c0;
  assign nS_st4_b51_c0 = nS_st3_b51_c0;
  assign nS_st4_b52_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b52_c0 : nS_st3_b52_c1;
  assign nS_st4_b53_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b53_c0 : nS_st3_b53_c1;
  assign nS_st4_b54_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b54_c0 : nS_st3_b54_c1;
  assign nS_st4_b55_c0 = (nC_st3_b51_c0 == 0) ? nS_st3_b55_c0 : nS_st3_b55_c1;
  assign nS_st4_b56_c0 = nS_st3_b56_c0;
  assign nS_st4_b57_c0 = nS_st3_b57_c0;
  assign nS_st4_b58_c0 = nS_st3_b58_c0;
  assign nS_st4_b59_c0 = nS_st3_b59_c0;
  assign nS_st4_b60_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b60_c0 : nS_st3_b60_c1;
  assign nS_st4_b61_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b61_c0 : nS_st3_b61_c1;
  assign nS_st4_b62_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b62_c0 : nS_st3_b62_c1;
  assign nS_st4_b63_c0 = (nC_st3_b59_c0 == 0) ? nS_st3_b63_c0 : nS_st3_b63_c1;
  assign nS_st4_b0_c1 = nS_st3_b0_c1;
  assign nS_st4_b1_c1 = nS_st3_b1_c1;
  assign nS_st4_b2_c1 = nS_st3_b2_c1;
  assign nS_st4_b3_c1 = nS_st3_b3_c1;
  assign nS_st4_b4_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b4_c0 : nS_st3_b4_c1;
  assign nS_st4_b5_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b5_c0 : nS_st3_b5_c1;
  assign nS_st4_b6_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b6_c0 : nS_st3_b6_c1;
  assign nS_st4_b7_c1 = (nC_st3_b3_c1 == 0) ? nS_st3_b7_c0 : nS_st3_b7_c1;
  assign nS_st4_b8_c1 = nS_st3_b8_c1;
  assign nS_st4_b9_c1 = nS_st3_b9_c1;
  assign nS_st4_b10_c1 = nS_st3_b10_c1;
  assign nS_st4_b11_c1 = nS_st3_b11_c1;
  assign nS_st4_b12_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b12_c0 : nS_st3_b12_c1;
  assign nS_st4_b13_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b13_c0 : nS_st3_b13_c1;
  assign nS_st4_b14_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b14_c0 : nS_st3_b14_c1;
  assign nS_st4_b15_c1 = (nC_st3_b11_c1 == 0) ? nS_st3_b15_c0 : nS_st3_b15_c1;
  assign nS_st4_b16_c1 = nS_st3_b16_c1;
  assign nS_st4_b17_c1 = nS_st3_b17_c1;
  assign nS_st4_b18_c1 = nS_st3_b18_c1;
  assign nS_st4_b19_c1 = nS_st3_b19_c1;
  assign nS_st4_b20_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b20_c0 : nS_st3_b20_c1;
  assign nS_st4_b21_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b21_c0 : nS_st3_b21_c1;
  assign nS_st4_b22_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b22_c0 : nS_st3_b22_c1;
  assign nS_st4_b23_c1 = (nC_st3_b19_c1 == 0) ? nS_st3_b23_c0 : nS_st3_b23_c1;
  assign nS_st4_b24_c1 = nS_st3_b24_c1;
  assign nS_st4_b25_c1 = nS_st3_b25_c1;
  assign nS_st4_b26_c1 = nS_st3_b26_c1;
  assign nS_st4_b27_c1 = nS_st3_b27_c1;
  assign nS_st4_b28_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b28_c0 : nS_st3_b28_c1;
  assign nS_st4_b29_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b29_c0 : nS_st3_b29_c1;
  assign nS_st4_b30_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b30_c0 : nS_st3_b30_c1;
  assign nS_st4_b31_c1 = (nC_st3_b27_c1 == 0) ? nS_st3_b31_c0 : nS_st3_b31_c1;
  assign nS_st4_b32_c1 = nS_st3_b32_c1;
  assign nS_st4_b33_c1 = nS_st3_b33_c1;
  assign nS_st4_b34_c1 = nS_st3_b34_c1;
  assign nS_st4_b35_c1 = nS_st3_b35_c1;
  assign nS_st4_b36_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b36_c0 : nS_st3_b36_c1;
  assign nS_st4_b37_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b37_c0 : nS_st3_b37_c1;
  assign nS_st4_b38_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b38_c0 : nS_st3_b38_c1;
  assign nS_st4_b39_c1 = (nC_st3_b35_c1 == 0) ? nS_st3_b39_c0 : nS_st3_b39_c1;
  assign nS_st4_b40_c1 = nS_st3_b40_c1;
  assign nS_st4_b41_c1 = nS_st3_b41_c1;
  assign nS_st4_b42_c1 = nS_st3_b42_c1;
  assign nS_st4_b43_c1 = nS_st3_b43_c1;
  assign nS_st4_b44_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b44_c0 : nS_st3_b44_c1;
  assign nS_st4_b45_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b45_c0 : nS_st3_b45_c1;
  assign nS_st4_b46_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b46_c0 : nS_st3_b46_c1;
  assign nS_st4_b47_c1 = (nC_st3_b43_c1 == 0) ? nS_st3_b47_c0 : nS_st3_b47_c1;
  assign nS_st4_b48_c1 = nS_st3_b48_c1;
  assign nS_st4_b49_c1 = nS_st3_b49_c1;
  assign nS_st4_b50_c1 = nS_st3_b50_c1;
  assign nS_st4_b51_c1 = nS_st3_b51_c1;
  assign nS_st4_b52_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b52_c0 : nS_st3_b52_c1;
  assign nS_st4_b53_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b53_c0 : nS_st3_b53_c1;
  assign nS_st4_b54_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b54_c0 : nS_st3_b54_c1;
  assign nS_st4_b55_c1 = (nC_st3_b51_c1 == 0) ? nS_st3_b55_c0 : nS_st3_b55_c1;
  assign nS_st4_b56_c1 = nS_st3_b56_c1;
  assign nS_st4_b57_c1 = nS_st3_b57_c1;
  assign nS_st4_b58_c1 = nS_st3_b58_c1;
  assign nS_st4_b59_c1 = nS_st3_b59_c1;
  assign nS_st4_b60_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b60_c0 : nS_st3_b60_c1;
  assign nS_st4_b61_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b61_c0 : nS_st3_b61_c1;
  assign nS_st4_b62_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b62_c0 : nS_st3_b62_c1;
  assign nS_st4_b63_c1 = (nC_st3_b59_c1 == 0) ? nS_st3_b63_c0 : nS_st3_b63_c1;
  assign nC_st4_b7_c0 = (nC_st3_b3_c0 == 0) ? nC_st3_b7_c0 : nC_st3_b7_c1;
  assign nC_st4_b15_c0 = (nC_st3_b11_c0 == 0) ? nC_st3_b15_c0 : nC_st3_b15_c1;
  assign nC_st4_b23_c0 = (nC_st3_b19_c0 == 0) ? nC_st3_b23_c0 : nC_st3_b23_c1;
  assign nC_st4_b31_c0 = (nC_st3_b27_c0 == 0) ? nC_st3_b31_c0 : nC_st3_b31_c1;
  assign nC_st4_b39_c0 = (nC_st3_b35_c0 == 0) ? nC_st3_b39_c0 : nC_st3_b39_c1;
  assign nC_st4_b47_c0 = (nC_st3_b43_c0 == 0) ? nC_st3_b47_c0 : nC_st3_b47_c1;
  assign nC_st4_b55_c0 = (nC_st3_b51_c0 == 0) ? nC_st3_b55_c0 : nC_st3_b55_c1;
  assign nC_st4_b63_c0 = (nC_st3_b59_c0 == 0) ? nC_st3_b63_c0 : nC_st3_b63_c1;
  assign nC_st4_b7_c1 = (nC_st3_b3_c1 == 0) ? nC_st3_b7_c0 : nC_st3_b7_c1;
  assign nC_st4_b15_c1 = (nC_st3_b11_c1 == 0) ? nC_st3_b15_c0 : nC_st3_b15_c1;
  assign nC_st4_b23_c1 = (nC_st3_b19_c1 == 0) ? nC_st3_b23_c0 : nC_st3_b23_c1;
  assign nC_st4_b31_c1 = (nC_st3_b27_c1 == 0) ? nC_st3_b31_c0 : nC_st3_b31_c1;
  assign nC_st4_b39_c1 = (nC_st3_b35_c1 == 0) ? nC_st3_b39_c0 : nC_st3_b39_c1;
  assign nC_st4_b47_c1 = (nC_st3_b43_c1 == 0) ? nC_st3_b47_c0 : nC_st3_b47_c1;
  assign nC_st4_b55_c1 = (nC_st3_b51_c1 == 0) ? nC_st3_b55_c0 : nC_st3_b55_c1;
  assign nC_st4_b63_c1 = (nC_st3_b59_c1 == 0) ? nC_st3_b63_c0 : nC_st3_b63_c1;

  assign nS_st5_b0_c0 = nS_st4_b0_c0;
  assign nS_st5_b1_c0 = nS_st4_b1_c0;
  assign nS_st5_b2_c0 = nS_st4_b2_c0;
  assign nS_st5_b3_c0 = nS_st4_b3_c0;
  assign nS_st5_b4_c0 = nS_st4_b4_c0;
  assign nS_st5_b5_c0 = nS_st4_b5_c0;
  assign nS_st5_b6_c0 = nS_st4_b6_c0;
  assign nS_st5_b7_c0 = nS_st4_b7_c0;
  assign nS_st5_b8_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b8_c0 : nS_st4_b8_c1;
  assign nS_st5_b9_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b9_c0 : nS_st4_b9_c1;
  assign nS_st5_b10_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b10_c0 : nS_st4_b10_c1;
  assign nS_st5_b11_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b11_c0 : nS_st4_b11_c1;
  assign nS_st5_b12_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b12_c0 : nS_st4_b12_c1;
  assign nS_st5_b13_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b13_c0 : nS_st4_b13_c1;
  assign nS_st5_b14_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b14_c0 : nS_st4_b14_c1;
  assign nS_st5_b15_c0 = (nC_st4_b7_c0 == 0) ? nS_st4_b15_c0 : nS_st4_b15_c1;
  assign nS_st5_b16_c0 = nS_st4_b16_c0;
  assign nS_st5_b17_c0 = nS_st4_b17_c0;
  assign nS_st5_b18_c0 = nS_st4_b18_c0;
  assign nS_st5_b19_c0 = nS_st4_b19_c0;
  assign nS_st5_b20_c0 = nS_st4_b20_c0;
  assign nS_st5_b21_c0 = nS_st4_b21_c0;
  assign nS_st5_b22_c0 = nS_st4_b22_c0;
  assign nS_st5_b23_c0 = nS_st4_b23_c0;
  assign nS_st5_b24_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b24_c0 : nS_st4_b24_c1;
  assign nS_st5_b25_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b25_c0 : nS_st4_b25_c1;
  assign nS_st5_b26_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b26_c0 : nS_st4_b26_c1;
  assign nS_st5_b27_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b27_c0 : nS_st4_b27_c1;
  assign nS_st5_b28_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b28_c0 : nS_st4_b28_c1;
  assign nS_st5_b29_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b29_c0 : nS_st4_b29_c1;
  assign nS_st5_b30_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b30_c0 : nS_st4_b30_c1;
  assign nS_st5_b31_c0 = (nC_st4_b23_c0 == 0) ? nS_st4_b31_c0 : nS_st4_b31_c1;
  assign nS_st5_b32_c0 = nS_st4_b32_c0;
  assign nS_st5_b33_c0 = nS_st4_b33_c0;
  assign nS_st5_b34_c0 = nS_st4_b34_c0;
  assign nS_st5_b35_c0 = nS_st4_b35_c0;
  assign nS_st5_b36_c0 = nS_st4_b36_c0;
  assign nS_st5_b37_c0 = nS_st4_b37_c0;
  assign nS_st5_b38_c0 = nS_st4_b38_c0;
  assign nS_st5_b39_c0 = nS_st4_b39_c0;
  assign nS_st5_b40_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b40_c0 : nS_st4_b40_c1;
  assign nS_st5_b41_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b41_c0 : nS_st4_b41_c1;
  assign nS_st5_b42_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b42_c0 : nS_st4_b42_c1;
  assign nS_st5_b43_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b43_c0 : nS_st4_b43_c1;
  assign nS_st5_b44_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b44_c0 : nS_st4_b44_c1;
  assign nS_st5_b45_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b45_c0 : nS_st4_b45_c1;
  assign nS_st5_b46_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b46_c0 : nS_st4_b46_c1;
  assign nS_st5_b47_c0 = (nC_st4_b39_c0 == 0) ? nS_st4_b47_c0 : nS_st4_b47_c1;
  assign nS_st5_b48_c0 = nS_st4_b48_c0;
  assign nS_st5_b49_c0 = nS_st4_b49_c0;
  assign nS_st5_b50_c0 = nS_st4_b50_c0;
  assign nS_st5_b51_c0 = nS_st4_b51_c0;
  assign nS_st5_b52_c0 = nS_st4_b52_c0;
  assign nS_st5_b53_c0 = nS_st4_b53_c0;
  assign nS_st5_b54_c0 = nS_st4_b54_c0;
  assign nS_st5_b55_c0 = nS_st4_b55_c0;
  assign nS_st5_b56_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b56_c0 : nS_st4_b56_c1;
  assign nS_st5_b57_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b57_c0 : nS_st4_b57_c1;
  assign nS_st5_b58_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b58_c0 : nS_st4_b58_c1;
  assign nS_st5_b59_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b59_c0 : nS_st4_b59_c1;
  assign nS_st5_b60_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b60_c0 : nS_st4_b60_c1;
  assign nS_st5_b61_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b61_c0 : nS_st4_b61_c1;
  assign nS_st5_b62_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b62_c0 : nS_st4_b62_c1;
  assign nS_st5_b63_c0 = (nC_st4_b55_c0 == 0) ? nS_st4_b63_c0 : nS_st4_b63_c1;
  assign nS_st5_b0_c1 = nS_st4_b0_c1;
  assign nS_st5_b1_c1 = nS_st4_b1_c1;
  assign nS_st5_b2_c1 = nS_st4_b2_c1;
  assign nS_st5_b3_c1 = nS_st4_b3_c1;
  assign nS_st5_b4_c1 = nS_st4_b4_c1;
  assign nS_st5_b5_c1 = nS_st4_b5_c1;
  assign nS_st5_b6_c1 = nS_st4_b6_c1;
  assign nS_st5_b7_c1 = nS_st4_b7_c1;
  assign nS_st5_b8_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b8_c0 : nS_st4_b8_c1;
  assign nS_st5_b9_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b9_c0 : nS_st4_b9_c1;
  assign nS_st5_b10_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b10_c0 : nS_st4_b10_c1;
  assign nS_st5_b11_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b11_c0 : nS_st4_b11_c1;
  assign nS_st5_b12_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b12_c0 : nS_st4_b12_c1;
  assign nS_st5_b13_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b13_c0 : nS_st4_b13_c1;
  assign nS_st5_b14_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b14_c0 : nS_st4_b14_c1;
  assign nS_st5_b15_c1 = (nC_st4_b7_c1 == 0) ? nS_st4_b15_c0 : nS_st4_b15_c1;
  assign nS_st5_b16_c1 = nS_st4_b16_c1;
  assign nS_st5_b17_c1 = nS_st4_b17_c1;
  assign nS_st5_b18_c1 = nS_st4_b18_c1;
  assign nS_st5_b19_c1 = nS_st4_b19_c1;
  assign nS_st5_b20_c1 = nS_st4_b20_c1;
  assign nS_st5_b21_c1 = nS_st4_b21_c1;
  assign nS_st5_b22_c1 = nS_st4_b22_c1;
  assign nS_st5_b23_c1 = nS_st4_b23_c1;
  assign nS_st5_b24_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b24_c0 : nS_st4_b24_c1;
  assign nS_st5_b25_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b25_c0 : nS_st4_b25_c1;
  assign nS_st5_b26_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b26_c0 : nS_st4_b26_c1;
  assign nS_st5_b27_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b27_c0 : nS_st4_b27_c1;
  assign nS_st5_b28_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b28_c0 : nS_st4_b28_c1;
  assign nS_st5_b29_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b29_c0 : nS_st4_b29_c1;
  assign nS_st5_b30_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b30_c0 : nS_st4_b30_c1;
  assign nS_st5_b31_c1 = (nC_st4_b23_c1 == 0) ? nS_st4_b31_c0 : nS_st4_b31_c1;
  assign nS_st5_b32_c1 = nS_st4_b32_c1;
  assign nS_st5_b33_c1 = nS_st4_b33_c1;
  assign nS_st5_b34_c1 = nS_st4_b34_c1;
  assign nS_st5_b35_c1 = nS_st4_b35_c1;
  assign nS_st5_b36_c1 = nS_st4_b36_c1;
  assign nS_st5_b37_c1 = nS_st4_b37_c1;
  assign nS_st5_b38_c1 = nS_st4_b38_c1;
  assign nS_st5_b39_c1 = nS_st4_b39_c1;
  assign nS_st5_b40_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b40_c0 : nS_st4_b40_c1;
  assign nS_st5_b41_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b41_c0 : nS_st4_b41_c1;
  assign nS_st5_b42_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b42_c0 : nS_st4_b42_c1;
  assign nS_st5_b43_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b43_c0 : nS_st4_b43_c1;
  assign nS_st5_b44_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b44_c0 : nS_st4_b44_c1;
  assign nS_st5_b45_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b45_c0 : nS_st4_b45_c1;
  assign nS_st5_b46_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b46_c0 : nS_st4_b46_c1;
  assign nS_st5_b47_c1 = (nC_st4_b39_c1 == 0) ? nS_st4_b47_c0 : nS_st4_b47_c1;
  assign nS_st5_b48_c1 = nS_st4_b48_c1;
  assign nS_st5_b49_c1 = nS_st4_b49_c1;
  assign nS_st5_b50_c1 = nS_st4_b50_c1;
  assign nS_st5_b51_c1 = nS_st4_b51_c1;
  assign nS_st5_b52_c1 = nS_st4_b52_c1;
  assign nS_st5_b53_c1 = nS_st4_b53_c1;
  assign nS_st5_b54_c1 = nS_st4_b54_c1;
  assign nS_st5_b55_c1 = nS_st4_b55_c1;
  assign nS_st5_b56_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b56_c0 : nS_st4_b56_c1;
  assign nS_st5_b57_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b57_c0 : nS_st4_b57_c1;
  assign nS_st5_b58_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b58_c0 : nS_st4_b58_c1;
  assign nS_st5_b59_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b59_c0 : nS_st4_b59_c1;
  assign nS_st5_b60_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b60_c0 : nS_st4_b60_c1;
  assign nS_st5_b61_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b61_c0 : nS_st4_b61_c1;
  assign nS_st5_b62_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b62_c0 : nS_st4_b62_c1;
  assign nS_st5_b63_c1 = (nC_st4_b55_c1 == 0) ? nS_st4_b63_c0 : nS_st4_b63_c1;
  assign nC_st5_b15_c0 = (nC_st4_b7_c0 == 0) ? nC_st4_b15_c0 : nC_st4_b15_c1;
  assign nC_st5_b31_c0 = (nC_st4_b23_c0 == 0) ? nC_st4_b31_c0 : nC_st4_b31_c1;
  assign nC_st5_b47_c0 = (nC_st4_b39_c0 == 0) ? nC_st4_b47_c0 : nC_st4_b47_c1;
  assign nC_st5_b63_c0 = (nC_st4_b55_c0 == 0) ? nC_st4_b63_c0 : nC_st4_b63_c1;
  assign nC_st5_b15_c1 = (nC_st4_b7_c1 == 0) ? nC_st4_b15_c0 : nC_st4_b15_c1;
  assign nC_st5_b31_c1 = (nC_st4_b23_c1 == 0) ? nC_st4_b31_c0 : nC_st4_b31_c1;
  assign nC_st5_b47_c1 = (nC_st4_b39_c1 == 0) ? nC_st4_b47_c0 : nC_st4_b47_c1;
  assign nC_st5_b63_c1 = (nC_st4_b55_c1 == 0) ? nC_st4_b63_c0 : nC_st4_b63_c1;

  assign nS_st6_b0_c0 = nS_st5_b0_c0;
  assign nS_st6_b1_c0 = nS_st5_b1_c0;
  assign nS_st6_b2_c0 = nS_st5_b2_c0;
  assign nS_st6_b3_c0 = nS_st5_b3_c0;
  assign nS_st6_b4_c0 = nS_st5_b4_c0;
  assign nS_st6_b5_c0 = nS_st5_b5_c0;
  assign nS_st6_b6_c0 = nS_st5_b6_c0;
  assign nS_st6_b7_c0 = nS_st5_b7_c0;
  assign nS_st6_b8_c0 = nS_st5_b8_c0;
  assign nS_st6_b9_c0 = nS_st5_b9_c0;
  assign nS_st6_b10_c0 = nS_st5_b10_c0;
  assign nS_st6_b11_c0 = nS_st5_b11_c0;
  assign nS_st6_b12_c0 = nS_st5_b12_c0;
  assign nS_st6_b13_c0 = nS_st5_b13_c0;
  assign nS_st6_b14_c0 = nS_st5_b14_c0;
  assign nS_st6_b15_c0 = nS_st5_b15_c0;
  assign nS_st6_b16_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b16_c0 : nS_st5_b16_c1;
  assign nS_st6_b17_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b17_c0 : nS_st5_b17_c1;
  assign nS_st6_b18_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b18_c0 : nS_st5_b18_c1;
  assign nS_st6_b19_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b19_c0 : nS_st5_b19_c1;
  assign nS_st6_b20_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b20_c0 : nS_st5_b20_c1;
  assign nS_st6_b21_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b21_c0 : nS_st5_b21_c1;
  assign nS_st6_b22_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b22_c0 : nS_st5_b22_c1;
  assign nS_st6_b23_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b23_c0 : nS_st5_b23_c1;
  assign nS_st6_b24_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b24_c0 : nS_st5_b24_c1;
  assign nS_st6_b25_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b25_c0 : nS_st5_b25_c1;
  assign nS_st6_b26_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b26_c0 : nS_st5_b26_c1;
  assign nS_st6_b27_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b27_c0 : nS_st5_b27_c1;
  assign nS_st6_b28_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b28_c0 : nS_st5_b28_c1;
  assign nS_st6_b29_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b29_c0 : nS_st5_b29_c1;
  assign nS_st6_b30_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b30_c0 : nS_st5_b30_c1;
  assign nS_st6_b31_c0 = (nC_st5_b15_c0 == 0) ? nS_st5_b31_c0 : nS_st5_b31_c1;
  assign nS_st6_b32_c0 = nS_st5_b32_c0;
  assign nS_st6_b33_c0 = nS_st5_b33_c0;
  assign nS_st6_b34_c0 = nS_st5_b34_c0;
  assign nS_st6_b35_c0 = nS_st5_b35_c0;
  assign nS_st6_b36_c0 = nS_st5_b36_c0;
  assign nS_st6_b37_c0 = nS_st5_b37_c0;
  assign nS_st6_b38_c0 = nS_st5_b38_c0;
  assign nS_st6_b39_c0 = nS_st5_b39_c0;
  assign nS_st6_b40_c0 = nS_st5_b40_c0;
  assign nS_st6_b41_c0 = nS_st5_b41_c0;
  assign nS_st6_b42_c0 = nS_st5_b42_c0;
  assign nS_st6_b43_c0 = nS_st5_b43_c0;
  assign nS_st6_b44_c0 = nS_st5_b44_c0;
  assign nS_st6_b45_c0 = nS_st5_b45_c0;
  assign nS_st6_b46_c0 = nS_st5_b46_c0;
  assign nS_st6_b47_c0 = nS_st5_b47_c0;
  assign nS_st6_b48_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b48_c0 : nS_st5_b48_c1;
  assign nS_st6_b49_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b49_c0 : nS_st5_b49_c1;
  assign nS_st6_b50_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b50_c0 : nS_st5_b50_c1;
  assign nS_st6_b51_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b51_c0 : nS_st5_b51_c1;
  assign nS_st6_b52_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b52_c0 : nS_st5_b52_c1;
  assign nS_st6_b53_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b53_c0 : nS_st5_b53_c1;
  assign nS_st6_b54_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b54_c0 : nS_st5_b54_c1;
  assign nS_st6_b55_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b55_c0 : nS_st5_b55_c1;
  assign nS_st6_b56_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b56_c0 : nS_st5_b56_c1;
  assign nS_st6_b57_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b57_c0 : nS_st5_b57_c1;
  assign nS_st6_b58_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b58_c0 : nS_st5_b58_c1;
  assign nS_st6_b59_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b59_c0 : nS_st5_b59_c1;
  assign nS_st6_b60_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b60_c0 : nS_st5_b60_c1;
  assign nS_st6_b61_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b61_c0 : nS_st5_b61_c1;
  assign nS_st6_b62_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b62_c0 : nS_st5_b62_c1;
  assign nS_st6_b63_c0 = (nC_st5_b47_c0 == 0) ? nS_st5_b63_c0 : nS_st5_b63_c1;
  assign nS_st6_b0_c1 = nS_st5_b0_c1;
  assign nS_st6_b1_c1 = nS_st5_b1_c1;
  assign nS_st6_b2_c1 = nS_st5_b2_c1;
  assign nS_st6_b3_c1 = nS_st5_b3_c1;
  assign nS_st6_b4_c1 = nS_st5_b4_c1;
  assign nS_st6_b5_c1 = nS_st5_b5_c1;
  assign nS_st6_b6_c1 = nS_st5_b6_c1;
  assign nS_st6_b7_c1 = nS_st5_b7_c1;
  assign nS_st6_b8_c1 = nS_st5_b8_c1;
  assign nS_st6_b9_c1 = nS_st5_b9_c1;
  assign nS_st6_b10_c1 = nS_st5_b10_c1;
  assign nS_st6_b11_c1 = nS_st5_b11_c1;
  assign nS_st6_b12_c1 = nS_st5_b12_c1;
  assign nS_st6_b13_c1 = nS_st5_b13_c1;
  assign nS_st6_b14_c1 = nS_st5_b14_c1;
  assign nS_st6_b15_c1 = nS_st5_b15_c1;
  assign nS_st6_b16_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b16_c0 : nS_st5_b16_c1;
  assign nS_st6_b17_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b17_c0 : nS_st5_b17_c1;
  assign nS_st6_b18_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b18_c0 : nS_st5_b18_c1;
  assign nS_st6_b19_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b19_c0 : nS_st5_b19_c1;
  assign nS_st6_b20_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b20_c0 : nS_st5_b20_c1;
  assign nS_st6_b21_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b21_c0 : nS_st5_b21_c1;
  assign nS_st6_b22_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b22_c0 : nS_st5_b22_c1;
  assign nS_st6_b23_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b23_c0 : nS_st5_b23_c1;
  assign nS_st6_b24_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b24_c0 : nS_st5_b24_c1;
  assign nS_st6_b25_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b25_c0 : nS_st5_b25_c1;
  assign nS_st6_b26_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b26_c0 : nS_st5_b26_c1;
  assign nS_st6_b27_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b27_c0 : nS_st5_b27_c1;
  assign nS_st6_b28_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b28_c0 : nS_st5_b28_c1;
  assign nS_st6_b29_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b29_c0 : nS_st5_b29_c1;
  assign nS_st6_b30_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b30_c0 : nS_st5_b30_c1;
  assign nS_st6_b31_c1 = (nC_st5_b15_c1 == 0) ? nS_st5_b31_c0 : nS_st5_b31_c1;
  assign nS_st6_b32_c1 = nS_st5_b32_c1;
  assign nS_st6_b33_c1 = nS_st5_b33_c1;
  assign nS_st6_b34_c1 = nS_st5_b34_c1;
  assign nS_st6_b35_c1 = nS_st5_b35_c1;
  assign nS_st6_b36_c1 = nS_st5_b36_c1;
  assign nS_st6_b37_c1 = nS_st5_b37_c1;
  assign nS_st6_b38_c1 = nS_st5_b38_c1;
  assign nS_st6_b39_c1 = nS_st5_b39_c1;
  assign nS_st6_b40_c1 = nS_st5_b40_c1;
  assign nS_st6_b41_c1 = nS_st5_b41_c1;
  assign nS_st6_b42_c1 = nS_st5_b42_c1;
  assign nS_st6_b43_c1 = nS_st5_b43_c1;
  assign nS_st6_b44_c1 = nS_st5_b44_c1;
  assign nS_st6_b45_c1 = nS_st5_b45_c1;
  assign nS_st6_b46_c1 = nS_st5_b46_c1;
  assign nS_st6_b47_c1 = nS_st5_b47_c1;
  assign nS_st6_b48_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b48_c0 : nS_st5_b48_c1;
  assign nS_st6_b49_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b49_c0 : nS_st5_b49_c1;
  assign nS_st6_b50_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b50_c0 : nS_st5_b50_c1;
  assign nS_st6_b51_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b51_c0 : nS_st5_b51_c1;
  assign nS_st6_b52_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b52_c0 : nS_st5_b52_c1;
  assign nS_st6_b53_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b53_c0 : nS_st5_b53_c1;
  assign nS_st6_b54_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b54_c0 : nS_st5_b54_c1;
  assign nS_st6_b55_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b55_c0 : nS_st5_b55_c1;
  assign nS_st6_b56_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b56_c0 : nS_st5_b56_c1;
  assign nS_st6_b57_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b57_c0 : nS_st5_b57_c1;
  assign nS_st6_b58_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b58_c0 : nS_st5_b58_c1;
  assign nS_st6_b59_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b59_c0 : nS_st5_b59_c1;
  assign nS_st6_b60_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b60_c0 : nS_st5_b60_c1;
  assign nS_st6_b61_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b61_c0 : nS_st5_b61_c1;
  assign nS_st6_b62_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b62_c0 : nS_st5_b62_c1;
  assign nS_st6_b63_c1 = (nC_st5_b47_c1 == 0) ? nS_st5_b63_c0 : nS_st5_b63_c1;
  assign nC_st6_b31_c0 = (nC_st5_b15_c0 == 0) ? nC_st5_b31_c0 : nC_st5_b31_c1;
  assign nC_st6_b63_c0 = (nC_st5_b47_c0 == 0) ? nC_st5_b63_c0 : nC_st5_b63_c1;
  assign nC_st6_b31_c1 = (nC_st5_b15_c1 == 0) ? nC_st5_b31_c0 : nC_st5_b31_c1;
  assign nC_st6_b63_c1 = (nC_st5_b47_c1 == 0) ? nC_st5_b63_c0 : nC_st5_b63_c1;

  assign nS_st7_b0_c0 = nS_st6_b0_c0;
  assign nS_st7_b1_c0 = nS_st6_b1_c0;
  assign nS_st7_b2_c0 = nS_st6_b2_c0;
  assign nS_st7_b3_c0 = nS_st6_b3_c0;
  assign nS_st7_b4_c0 = nS_st6_b4_c0;
  assign nS_st7_b5_c0 = nS_st6_b5_c0;
  assign nS_st7_b6_c0 = nS_st6_b6_c0;
  assign nS_st7_b7_c0 = nS_st6_b7_c0;
  assign nS_st7_b8_c0 = nS_st6_b8_c0;
  assign nS_st7_b9_c0 = nS_st6_b9_c0;
  assign nS_st7_b10_c0 = nS_st6_b10_c0;
  assign nS_st7_b11_c0 = nS_st6_b11_c0;
  assign nS_st7_b12_c0 = nS_st6_b12_c0;
  assign nS_st7_b13_c0 = nS_st6_b13_c0;
  assign nS_st7_b14_c0 = nS_st6_b14_c0;
  assign nS_st7_b15_c0 = nS_st6_b15_c0;
  assign nS_st7_b16_c0 = nS_st6_b16_c0;
  assign nS_st7_b17_c0 = nS_st6_b17_c0;
  assign nS_st7_b18_c0 = nS_st6_b18_c0;
  assign nS_st7_b19_c0 = nS_st6_b19_c0;
  assign nS_st7_b20_c0 = nS_st6_b20_c0;
  assign nS_st7_b21_c0 = nS_st6_b21_c0;
  assign nS_st7_b22_c0 = nS_st6_b22_c0;
  assign nS_st7_b23_c0 = nS_st6_b23_c0;
  assign nS_st7_b24_c0 = nS_st6_b24_c0;
  assign nS_st7_b25_c0 = nS_st6_b25_c0;
  assign nS_st7_b26_c0 = nS_st6_b26_c0;
  assign nS_st7_b27_c0 = nS_st6_b27_c0;
  assign nS_st7_b28_c0 = nS_st6_b28_c0;
  assign nS_st7_b29_c0 = nS_st6_b29_c0;
  assign nS_st7_b30_c0 = nS_st6_b30_c0;
  assign nS_st7_b31_c0 = nS_st6_b31_c0;
  assign nS_st7_b32_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b32_c0 : nS_st6_b32_c1;
  assign nS_st7_b33_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b33_c0 : nS_st6_b33_c1;
  assign nS_st7_b34_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b34_c0 : nS_st6_b34_c1;
  assign nS_st7_b35_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b35_c0 : nS_st6_b35_c1;
  assign nS_st7_b36_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b36_c0 : nS_st6_b36_c1;
  assign nS_st7_b37_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b37_c0 : nS_st6_b37_c1;
  assign nS_st7_b38_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b38_c0 : nS_st6_b38_c1;
  assign nS_st7_b39_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b39_c0 : nS_st6_b39_c1;
  assign nS_st7_b40_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b40_c0 : nS_st6_b40_c1;
  assign nS_st7_b41_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b41_c0 : nS_st6_b41_c1;
  assign nS_st7_b42_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b42_c0 : nS_st6_b42_c1;
  assign nS_st7_b43_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b43_c0 : nS_st6_b43_c1;
  assign nS_st7_b44_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b44_c0 : nS_st6_b44_c1;
  assign nS_st7_b45_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b45_c0 : nS_st6_b45_c1;
  assign nS_st7_b46_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b46_c0 : nS_st6_b46_c1;
  assign nS_st7_b47_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b47_c0 : nS_st6_b47_c1;
  assign nS_st7_b48_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b48_c0 : nS_st6_b48_c1;
  assign nS_st7_b49_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b49_c0 : nS_st6_b49_c1;
  assign nS_st7_b50_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b50_c0 : nS_st6_b50_c1;
  assign nS_st7_b51_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b51_c0 : nS_st6_b51_c1;
  assign nS_st7_b52_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b52_c0 : nS_st6_b52_c1;
  assign nS_st7_b53_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b53_c0 : nS_st6_b53_c1;
  assign nS_st7_b54_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b54_c0 : nS_st6_b54_c1;
  assign nS_st7_b55_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b55_c0 : nS_st6_b55_c1;
  assign nS_st7_b56_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b56_c0 : nS_st6_b56_c1;
  assign nS_st7_b57_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b57_c0 : nS_st6_b57_c1;
  assign nS_st7_b58_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b58_c0 : nS_st6_b58_c1;
  assign nS_st7_b59_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b59_c0 : nS_st6_b59_c1;
  assign nS_st7_b60_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b60_c0 : nS_st6_b60_c1;
  assign nS_st7_b61_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b61_c0 : nS_st6_b61_c1;
  assign nS_st7_b62_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b62_c0 : nS_st6_b62_c1;
  assign nS_st7_b63_c0 = (nC_st6_b31_c0 == 0) ? nS_st6_b63_c0 : nS_st6_b63_c1;
  assign nS_st7_b0_c1 = nS_st6_b0_c1;
  assign nS_st7_b1_c1 = nS_st6_b1_c1;
  assign nS_st7_b2_c1 = nS_st6_b2_c1;
  assign nS_st7_b3_c1 = nS_st6_b3_c1;
  assign nS_st7_b4_c1 = nS_st6_b4_c1;
  assign nS_st7_b5_c1 = nS_st6_b5_c1;
  assign nS_st7_b6_c1 = nS_st6_b6_c1;
  assign nS_st7_b7_c1 = nS_st6_b7_c1;
  assign nS_st7_b8_c1 = nS_st6_b8_c1;
  assign nS_st7_b9_c1 = nS_st6_b9_c1;
  assign nS_st7_b10_c1 = nS_st6_b10_c1;
  assign nS_st7_b11_c1 = nS_st6_b11_c1;
  assign nS_st7_b12_c1 = nS_st6_b12_c1;
  assign nS_st7_b13_c1 = nS_st6_b13_c1;
  assign nS_st7_b14_c1 = nS_st6_b14_c1;
  assign nS_st7_b15_c1 = nS_st6_b15_c1;
  assign nS_st7_b16_c1 = nS_st6_b16_c1;
  assign nS_st7_b17_c1 = nS_st6_b17_c1;
  assign nS_st7_b18_c1 = nS_st6_b18_c1;
  assign nS_st7_b19_c1 = nS_st6_b19_c1;
  assign nS_st7_b20_c1 = nS_st6_b20_c1;
  assign nS_st7_b21_c1 = nS_st6_b21_c1;
  assign nS_st7_b22_c1 = nS_st6_b22_c1;
  assign nS_st7_b23_c1 = nS_st6_b23_c1;
  assign nS_st7_b24_c1 = nS_st6_b24_c1;
  assign nS_st7_b25_c1 = nS_st6_b25_c1;
  assign nS_st7_b26_c1 = nS_st6_b26_c1;
  assign nS_st7_b27_c1 = nS_st6_b27_c1;
  assign nS_st7_b28_c1 = nS_st6_b28_c1;
  assign nS_st7_b29_c1 = nS_st6_b29_c1;
  assign nS_st7_b30_c1 = nS_st6_b30_c1;
  assign nS_st7_b31_c1 = nS_st6_b31_c1;
  assign nS_st7_b32_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b32_c0 : nS_st6_b32_c1;
  assign nS_st7_b33_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b33_c0 : nS_st6_b33_c1;
  assign nS_st7_b34_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b34_c0 : nS_st6_b34_c1;
  assign nS_st7_b35_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b35_c0 : nS_st6_b35_c1;
  assign nS_st7_b36_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b36_c0 : nS_st6_b36_c1;
  assign nS_st7_b37_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b37_c0 : nS_st6_b37_c1;
  assign nS_st7_b38_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b38_c0 : nS_st6_b38_c1;
  assign nS_st7_b39_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b39_c0 : nS_st6_b39_c1;
  assign nS_st7_b40_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b40_c0 : nS_st6_b40_c1;
  assign nS_st7_b41_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b41_c0 : nS_st6_b41_c1;
  assign nS_st7_b42_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b42_c0 : nS_st6_b42_c1;
  assign nS_st7_b43_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b43_c0 : nS_st6_b43_c1;
  assign nS_st7_b44_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b44_c0 : nS_st6_b44_c1;
  assign nS_st7_b45_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b45_c0 : nS_st6_b45_c1;
  assign nS_st7_b46_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b46_c0 : nS_st6_b46_c1;
  assign nS_st7_b47_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b47_c0 : nS_st6_b47_c1;
  assign nS_st7_b48_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b48_c0 : nS_st6_b48_c1;
  assign nS_st7_b49_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b49_c0 : nS_st6_b49_c1;
  assign nS_st7_b50_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b50_c0 : nS_st6_b50_c1;
  assign nS_st7_b51_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b51_c0 : nS_st6_b51_c1;
  assign nS_st7_b52_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b52_c0 : nS_st6_b52_c1;
  assign nS_st7_b53_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b53_c0 : nS_st6_b53_c1;
  assign nS_st7_b54_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b54_c0 : nS_st6_b54_c1;
  assign nS_st7_b55_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b55_c0 : nS_st6_b55_c1;
  assign nS_st7_b56_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b56_c0 : nS_st6_b56_c1;
  assign nS_st7_b57_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b57_c0 : nS_st6_b57_c1;
  assign nS_st7_b58_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b58_c0 : nS_st6_b58_c1;
  assign nS_st7_b59_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b59_c0 : nS_st6_b59_c1;
  assign nS_st7_b60_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b60_c0 : nS_st6_b60_c1;
  assign nS_st7_b61_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b61_c0 : nS_st6_b61_c1;
  assign nS_st7_b62_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b62_c0 : nS_st6_b62_c1;
  assign nS_st7_b63_c1 = (nC_st6_b31_c1 == 0) ? nS_st6_b63_c0 : nS_st6_b63_c1;
  assign nC_st7_b63_c0 = (nC_st6_b31_c0 == 0) ? nC_st6_b63_c0 : nC_st6_b63_c1;
  assign nC_st7_b63_c1 = (nC_st6_b31_c1 == 0) ? nC_st6_b63_c0 : nC_st6_b63_c1;

  assign out_S[0] = (in_CI == 0) ? nS_st7_b0_c0 : nS_st7_b0_c1;
  assign out_S[1] = (in_CI == 0) ? nS_st7_b1_c0 : nS_st7_b1_c1;
  assign out_S[2] = (in_CI == 0) ? nS_st7_b2_c0 : nS_st7_b2_c1;
  assign out_S[3] = (in_CI == 0) ? nS_st7_b3_c0 : nS_st7_b3_c1;
  assign out_S[4] = (in_CI == 0) ? nS_st7_b4_c0 : nS_st7_b4_c1;
  assign out_S[5] = (in_CI == 0) ? nS_st7_b5_c0 : nS_st7_b5_c1;
  assign out_S[6] = (in_CI == 0) ? nS_st7_b6_c0 : nS_st7_b6_c1;
  assign out_S[7] = (in_CI == 0) ? nS_st7_b7_c0 : nS_st7_b7_c1;
  assign out_S[8] = (in_CI == 0) ? nS_st7_b8_c0 : nS_st7_b8_c1;
  assign out_S[9] = (in_CI == 0) ? nS_st7_b9_c0 : nS_st7_b9_c1;
  assign out_S[10] = (in_CI == 0) ? nS_st7_b10_c0 : nS_st7_b10_c1;
  assign out_S[11] = (in_CI == 0) ? nS_st7_b11_c0 : nS_st7_b11_c1;
  assign out_S[12] = (in_CI == 0) ? nS_st7_b12_c0 : nS_st7_b12_c1;
  assign out_S[13] = (in_CI == 0) ? nS_st7_b13_c0 : nS_st7_b13_c1;
  assign out_S[14] = (in_CI == 0) ? nS_st7_b14_c0 : nS_st7_b14_c1;
  assign out_S[15] = (in_CI == 0) ? nS_st7_b15_c0 : nS_st7_b15_c1;
  assign out_S[16] = (in_CI == 0) ? nS_st7_b16_c0 : nS_st7_b16_c1;
  assign out_S[17] = (in_CI == 0) ? nS_st7_b17_c0 : nS_st7_b17_c1;
  assign out_S[18] = (in_CI == 0) ? nS_st7_b18_c0 : nS_st7_b18_c1;
  assign out_S[19] = (in_CI == 0) ? nS_st7_b19_c0 : nS_st7_b19_c1;
  assign out_S[20] = (in_CI == 0) ? nS_st7_b20_c0 : nS_st7_b20_c1;
  assign out_S[21] = (in_CI == 0) ? nS_st7_b21_c0 : nS_st7_b21_c1;
  assign out_S[22] = (in_CI == 0) ? nS_st7_b22_c0 : nS_st7_b22_c1;
  assign out_S[23] = (in_CI == 0) ? nS_st7_b23_c0 : nS_st7_b23_c1;
  assign out_S[24] = (in_CI == 0) ? nS_st7_b24_c0 : nS_st7_b24_c1;
  assign out_S[25] = (in_CI == 0) ? nS_st7_b25_c0 : nS_st7_b25_c1;
  assign out_S[26] = (in_CI == 0) ? nS_st7_b26_c0 : nS_st7_b26_c1;
  assign out_S[27] = (in_CI == 0) ? nS_st7_b27_c0 : nS_st7_b27_c1;
  assign out_S[28] = (in_CI == 0) ? nS_st7_b28_c0 : nS_st7_b28_c1;
  assign out_S[29] = (in_CI == 0) ? nS_st7_b29_c0 : nS_st7_b29_c1;
  assign out_S[30] = (in_CI == 0) ? nS_st7_b30_c0 : nS_st7_b30_c1;
  assign out_S[31] = (in_CI == 0) ? nS_st7_b31_c0 : nS_st7_b31_c1;
  assign out_S[32] = (in_CI == 0) ? nS_st7_b32_c0 : nS_st7_b32_c1;
  assign out_S[33] = (in_CI == 0) ? nS_st7_b33_c0 : nS_st7_b33_c1;
  assign out_S[34] = (in_CI == 0) ? nS_st7_b34_c0 : nS_st7_b34_c1;
  assign out_S[35] = (in_CI == 0) ? nS_st7_b35_c0 : nS_st7_b35_c1;
  assign out_S[36] = (in_CI == 0) ? nS_st7_b36_c0 : nS_st7_b36_c1;
  assign out_S[37] = (in_CI == 0) ? nS_st7_b37_c0 : nS_st7_b37_c1;
  assign out_S[38] = (in_CI == 0) ? nS_st7_b38_c0 : nS_st7_b38_c1;
  assign out_S[39] = (in_CI == 0) ? nS_st7_b39_c0 : nS_st7_b39_c1;
  assign out_S[40] = (in_CI == 0) ? nS_st7_b40_c0 : nS_st7_b40_c1;
  assign out_S[41] = (in_CI == 0) ? nS_st7_b41_c0 : nS_st7_b41_c1;
  assign out_S[42] = (in_CI == 0) ? nS_st7_b42_c0 : nS_st7_b42_c1;
  assign out_S[43] = (in_CI == 0) ? nS_st7_b43_c0 : nS_st7_b43_c1;
  assign out_S[44] = (in_CI == 0) ? nS_st7_b44_c0 : nS_st7_b44_c1;
  assign out_S[45] = (in_CI == 0) ? nS_st7_b45_c0 : nS_st7_b45_c1;
  assign out_S[46] = (in_CI == 0) ? nS_st7_b46_c0 : nS_st7_b46_c1;
  assign out_S[47] = (in_CI == 0) ? nS_st7_b47_c0 : nS_st7_b47_c1;
  assign out_S[48] = (in_CI == 0) ? nS_st7_b48_c0 : nS_st7_b48_c1;
  assign out_S[49] = (in_CI == 0) ? nS_st7_b49_c0 : nS_st7_b49_c1;
  assign out_S[50] = (in_CI == 0) ? nS_st7_b50_c0 : nS_st7_b50_c1;
  assign out_S[51] = (in_CI == 0) ? nS_st7_b51_c0 : nS_st7_b51_c1;
  assign out_S[52] = (in_CI == 0) ? nS_st7_b52_c0 : nS_st7_b52_c1;
  assign out_S[53] = (in_CI == 0) ? nS_st7_b53_c0 : nS_st7_b53_c1;
  assign out_S[54] = (in_CI == 0) ? nS_st7_b54_c0 : nS_st7_b54_c1;
  assign out_S[55] = (in_CI == 0) ? nS_st7_b55_c0 : nS_st7_b55_c1;
  assign out_S[56] = (in_CI == 0) ? nS_st7_b56_c0 : nS_st7_b56_c1;
  assign out_S[57] = (in_CI == 0) ? nS_st7_b57_c0 : nS_st7_b57_c1;
  assign out_S[58] = (in_CI == 0) ? nS_st7_b58_c0 : nS_st7_b58_c1;
  assign out_S[59] = (in_CI == 0) ? nS_st7_b59_c0 : nS_st7_b59_c1;
  assign out_S[60] = (in_CI == 0) ? nS_st7_b60_c0 : nS_st7_b60_c1;
  assign out_S[61] = (in_CI == 0) ? nS_st7_b61_c0 : nS_st7_b61_c1;
  assign out_S[62] = (in_CI == 0) ? nS_st7_b62_c0 : nS_st7_b62_c1;
  assign out_S[63] = (in_CI == 0) ? nS_st7_b63_c0 : nS_st7_b63_c1;
  assign out_CO = (in_CI == 0) ? nC_st7_b63_c0 : nC_st7_b63_c1;
endmodule

