module VKSA_256 (in_A, in_B, in_CI, out_S, out_CO);
  input [255:0] in_A, in_B;
  input in_CI;
  output [255:0] out_S;
  output out_CO;

  assign nG_0_0 = in_A[0] & in_B[0];
  assign nP_0_0 = in_A[0] ^ in_B[0];
  assign nG_1_1 = in_A[1] & in_B[1];
  assign nP_1_1 = in_A[1] ^ in_B[1];
  assign nG_2_2 = in_A[2] & in_B[2];
  assign nP_2_2 = in_A[2] ^ in_B[2];
  assign nG_3_3 = in_A[3] & in_B[3];
  assign nP_3_3 = in_A[3] ^ in_B[3];
  assign nG_4_4 = in_A[4] & in_B[4];
  assign nP_4_4 = in_A[4] ^ in_B[4];
  assign nG_5_5 = in_A[5] & in_B[5];
  assign nP_5_5 = in_A[5] ^ in_B[5];
  assign nG_6_6 = in_A[6] & in_B[6];
  assign nP_6_6 = in_A[6] ^ in_B[6];
  assign nG_7_7 = in_A[7] & in_B[7];
  assign nP_7_7 = in_A[7] ^ in_B[7];
  assign nG_8_8 = in_A[8] & in_B[8];
  assign nP_8_8 = in_A[8] ^ in_B[8];
  assign nG_9_9 = in_A[9] & in_B[9];
  assign nP_9_9 = in_A[9] ^ in_B[9];
  assign nG_10_10 = in_A[10] & in_B[10];
  assign nP_10_10 = in_A[10] ^ in_B[10];
  assign nG_11_11 = in_A[11] & in_B[11];
  assign nP_11_11 = in_A[11] ^ in_B[11];
  assign nG_12_12 = in_A[12] & in_B[12];
  assign nP_12_12 = in_A[12] ^ in_B[12];
  assign nG_13_13 = in_A[13] & in_B[13];
  assign nP_13_13 = in_A[13] ^ in_B[13];
  assign nG_14_14 = in_A[14] & in_B[14];
  assign nP_14_14 = in_A[14] ^ in_B[14];
  assign nG_15_15 = in_A[15] & in_B[15];
  assign nP_15_15 = in_A[15] ^ in_B[15];
  assign nG_16_16 = in_A[16] & in_B[16];
  assign nP_16_16 = in_A[16] ^ in_B[16];
  assign nG_17_17 = in_A[17] & in_B[17];
  assign nP_17_17 = in_A[17] ^ in_B[17];
  assign nG_18_18 = in_A[18] & in_B[18];
  assign nP_18_18 = in_A[18] ^ in_B[18];
  assign nG_19_19 = in_A[19] & in_B[19];
  assign nP_19_19 = in_A[19] ^ in_B[19];
  assign nG_20_20 = in_A[20] & in_B[20];
  assign nP_20_20 = in_A[20] ^ in_B[20];
  assign nG_21_21 = in_A[21] & in_B[21];
  assign nP_21_21 = in_A[21] ^ in_B[21];
  assign nG_22_22 = in_A[22] & in_B[22];
  assign nP_22_22 = in_A[22] ^ in_B[22];
  assign nG_23_23 = in_A[23] & in_B[23];
  assign nP_23_23 = in_A[23] ^ in_B[23];
  assign nG_24_24 = in_A[24] & in_B[24];
  assign nP_24_24 = in_A[24] ^ in_B[24];
  assign nG_25_25 = in_A[25] & in_B[25];
  assign nP_25_25 = in_A[25] ^ in_B[25];
  assign nG_26_26 = in_A[26] & in_B[26];
  assign nP_26_26 = in_A[26] ^ in_B[26];
  assign nG_27_27 = in_A[27] & in_B[27];
  assign nP_27_27 = in_A[27] ^ in_B[27];
  assign nG_28_28 = in_A[28] & in_B[28];
  assign nP_28_28 = in_A[28] ^ in_B[28];
  assign nG_29_29 = in_A[29] & in_B[29];
  assign nP_29_29 = in_A[29] ^ in_B[29];
  assign nG_30_30 = in_A[30] & in_B[30];
  assign nP_30_30 = in_A[30] ^ in_B[30];
  assign nG_31_31 = in_A[31] & in_B[31];
  assign nP_31_31 = in_A[31] ^ in_B[31];
  assign nG_32_32 = in_A[32] & in_B[32];
  assign nP_32_32 = in_A[32] ^ in_B[32];
  assign nG_33_33 = in_A[33] & in_B[33];
  assign nP_33_33 = in_A[33] ^ in_B[33];
  assign nG_34_34 = in_A[34] & in_B[34];
  assign nP_34_34 = in_A[34] ^ in_B[34];
  assign nG_35_35 = in_A[35] & in_B[35];
  assign nP_35_35 = in_A[35] ^ in_B[35];
  assign nG_36_36 = in_A[36] & in_B[36];
  assign nP_36_36 = in_A[36] ^ in_B[36];
  assign nG_37_37 = in_A[37] & in_B[37];
  assign nP_37_37 = in_A[37] ^ in_B[37];
  assign nG_38_38 = in_A[38] & in_B[38];
  assign nP_38_38 = in_A[38] ^ in_B[38];
  assign nG_39_39 = in_A[39] & in_B[39];
  assign nP_39_39 = in_A[39] ^ in_B[39];
  assign nG_40_40 = in_A[40] & in_B[40];
  assign nP_40_40 = in_A[40] ^ in_B[40];
  assign nG_41_41 = in_A[41] & in_B[41];
  assign nP_41_41 = in_A[41] ^ in_B[41];
  assign nG_42_42 = in_A[42] & in_B[42];
  assign nP_42_42 = in_A[42] ^ in_B[42];
  assign nG_43_43 = in_A[43] & in_B[43];
  assign nP_43_43 = in_A[43] ^ in_B[43];
  assign nG_44_44 = in_A[44] & in_B[44];
  assign nP_44_44 = in_A[44] ^ in_B[44];
  assign nG_45_45 = in_A[45] & in_B[45];
  assign nP_45_45 = in_A[45] ^ in_B[45];
  assign nG_46_46 = in_A[46] & in_B[46];
  assign nP_46_46 = in_A[46] ^ in_B[46];
  assign nG_47_47 = in_A[47] & in_B[47];
  assign nP_47_47 = in_A[47] ^ in_B[47];
  assign nG_48_48 = in_A[48] & in_B[48];
  assign nP_48_48 = in_A[48] ^ in_B[48];
  assign nG_49_49 = in_A[49] & in_B[49];
  assign nP_49_49 = in_A[49] ^ in_B[49];
  assign nG_50_50 = in_A[50] & in_B[50];
  assign nP_50_50 = in_A[50] ^ in_B[50];
  assign nG_51_51 = in_A[51] & in_B[51];
  assign nP_51_51 = in_A[51] ^ in_B[51];
  assign nG_52_52 = in_A[52] & in_B[52];
  assign nP_52_52 = in_A[52] ^ in_B[52];
  assign nG_53_53 = in_A[53] & in_B[53];
  assign nP_53_53 = in_A[53] ^ in_B[53];
  assign nG_54_54 = in_A[54] & in_B[54];
  assign nP_54_54 = in_A[54] ^ in_B[54];
  assign nG_55_55 = in_A[55] & in_B[55];
  assign nP_55_55 = in_A[55] ^ in_B[55];
  assign nG_56_56 = in_A[56] & in_B[56];
  assign nP_56_56 = in_A[56] ^ in_B[56];
  assign nG_57_57 = in_A[57] & in_B[57];
  assign nP_57_57 = in_A[57] ^ in_B[57];
  assign nG_58_58 = in_A[58] & in_B[58];
  assign nP_58_58 = in_A[58] ^ in_B[58];
  assign nG_59_59 = in_A[59] & in_B[59];
  assign nP_59_59 = in_A[59] ^ in_B[59];
  assign nG_60_60 = in_A[60] & in_B[60];
  assign nP_60_60 = in_A[60] ^ in_B[60];
  assign nG_61_61 = in_A[61] & in_B[61];
  assign nP_61_61 = in_A[61] ^ in_B[61];
  assign nG_62_62 = in_A[62] & in_B[62];
  assign nP_62_62 = in_A[62] ^ in_B[62];
  assign nG_63_63 = in_A[63] & in_B[63];
  assign nP_63_63 = in_A[63] ^ in_B[63];
  assign nG_64_64 = in_A[64] & in_B[64];
  assign nP_64_64 = in_A[64] ^ in_B[64];
  assign nG_65_65 = in_A[65] & in_B[65];
  assign nP_65_65 = in_A[65] ^ in_B[65];
  assign nG_66_66 = in_A[66] & in_B[66];
  assign nP_66_66 = in_A[66] ^ in_B[66];
  assign nG_67_67 = in_A[67] & in_B[67];
  assign nP_67_67 = in_A[67] ^ in_B[67];
  assign nG_68_68 = in_A[68] & in_B[68];
  assign nP_68_68 = in_A[68] ^ in_B[68];
  assign nG_69_69 = in_A[69] & in_B[69];
  assign nP_69_69 = in_A[69] ^ in_B[69];
  assign nG_70_70 = in_A[70] & in_B[70];
  assign nP_70_70 = in_A[70] ^ in_B[70];
  assign nG_71_71 = in_A[71] & in_B[71];
  assign nP_71_71 = in_A[71] ^ in_B[71];
  assign nG_72_72 = in_A[72] & in_B[72];
  assign nP_72_72 = in_A[72] ^ in_B[72];
  assign nG_73_73 = in_A[73] & in_B[73];
  assign nP_73_73 = in_A[73] ^ in_B[73];
  assign nG_74_74 = in_A[74] & in_B[74];
  assign nP_74_74 = in_A[74] ^ in_B[74];
  assign nG_75_75 = in_A[75] & in_B[75];
  assign nP_75_75 = in_A[75] ^ in_B[75];
  assign nG_76_76 = in_A[76] & in_B[76];
  assign nP_76_76 = in_A[76] ^ in_B[76];
  assign nG_77_77 = in_A[77] & in_B[77];
  assign nP_77_77 = in_A[77] ^ in_B[77];
  assign nG_78_78 = in_A[78] & in_B[78];
  assign nP_78_78 = in_A[78] ^ in_B[78];
  assign nG_79_79 = in_A[79] & in_B[79];
  assign nP_79_79 = in_A[79] ^ in_B[79];
  assign nG_80_80 = in_A[80] & in_B[80];
  assign nP_80_80 = in_A[80] ^ in_B[80];
  assign nG_81_81 = in_A[81] & in_B[81];
  assign nP_81_81 = in_A[81] ^ in_B[81];
  assign nG_82_82 = in_A[82] & in_B[82];
  assign nP_82_82 = in_A[82] ^ in_B[82];
  assign nG_83_83 = in_A[83] & in_B[83];
  assign nP_83_83 = in_A[83] ^ in_B[83];
  assign nG_84_84 = in_A[84] & in_B[84];
  assign nP_84_84 = in_A[84] ^ in_B[84];
  assign nG_85_85 = in_A[85] & in_B[85];
  assign nP_85_85 = in_A[85] ^ in_B[85];
  assign nG_86_86 = in_A[86] & in_B[86];
  assign nP_86_86 = in_A[86] ^ in_B[86];
  assign nG_87_87 = in_A[87] & in_B[87];
  assign nP_87_87 = in_A[87] ^ in_B[87];
  assign nG_88_88 = in_A[88] & in_B[88];
  assign nP_88_88 = in_A[88] ^ in_B[88];
  assign nG_89_89 = in_A[89] & in_B[89];
  assign nP_89_89 = in_A[89] ^ in_B[89];
  assign nG_90_90 = in_A[90] & in_B[90];
  assign nP_90_90 = in_A[90] ^ in_B[90];
  assign nG_91_91 = in_A[91] & in_B[91];
  assign nP_91_91 = in_A[91] ^ in_B[91];
  assign nG_92_92 = in_A[92] & in_B[92];
  assign nP_92_92 = in_A[92] ^ in_B[92];
  assign nG_93_93 = in_A[93] & in_B[93];
  assign nP_93_93 = in_A[93] ^ in_B[93];
  assign nG_94_94 = in_A[94] & in_B[94];
  assign nP_94_94 = in_A[94] ^ in_B[94];
  assign nG_95_95 = in_A[95] & in_B[95];
  assign nP_95_95 = in_A[95] ^ in_B[95];
  assign nG_96_96 = in_A[96] & in_B[96];
  assign nP_96_96 = in_A[96] ^ in_B[96];
  assign nG_97_97 = in_A[97] & in_B[97];
  assign nP_97_97 = in_A[97] ^ in_B[97];
  assign nG_98_98 = in_A[98] & in_B[98];
  assign nP_98_98 = in_A[98] ^ in_B[98];
  assign nG_99_99 = in_A[99] & in_B[99];
  assign nP_99_99 = in_A[99] ^ in_B[99];
  assign nG_100_100 = in_A[100] & in_B[100];
  assign nP_100_100 = in_A[100] ^ in_B[100];
  assign nG_101_101 = in_A[101] & in_B[101];
  assign nP_101_101 = in_A[101] ^ in_B[101];
  assign nG_102_102 = in_A[102] & in_B[102];
  assign nP_102_102 = in_A[102] ^ in_B[102];
  assign nG_103_103 = in_A[103] & in_B[103];
  assign nP_103_103 = in_A[103] ^ in_B[103];
  assign nG_104_104 = in_A[104] & in_B[104];
  assign nP_104_104 = in_A[104] ^ in_B[104];
  assign nG_105_105 = in_A[105] & in_B[105];
  assign nP_105_105 = in_A[105] ^ in_B[105];
  assign nG_106_106 = in_A[106] & in_B[106];
  assign nP_106_106 = in_A[106] ^ in_B[106];
  assign nG_107_107 = in_A[107] & in_B[107];
  assign nP_107_107 = in_A[107] ^ in_B[107];
  assign nG_108_108 = in_A[108] & in_B[108];
  assign nP_108_108 = in_A[108] ^ in_B[108];
  assign nG_109_109 = in_A[109] & in_B[109];
  assign nP_109_109 = in_A[109] ^ in_B[109];
  assign nG_110_110 = in_A[110] & in_B[110];
  assign nP_110_110 = in_A[110] ^ in_B[110];
  assign nG_111_111 = in_A[111] & in_B[111];
  assign nP_111_111 = in_A[111] ^ in_B[111];
  assign nG_112_112 = in_A[112] & in_B[112];
  assign nP_112_112 = in_A[112] ^ in_B[112];
  assign nG_113_113 = in_A[113] & in_B[113];
  assign nP_113_113 = in_A[113] ^ in_B[113];
  assign nG_114_114 = in_A[114] & in_B[114];
  assign nP_114_114 = in_A[114] ^ in_B[114];
  assign nG_115_115 = in_A[115] & in_B[115];
  assign nP_115_115 = in_A[115] ^ in_B[115];
  assign nG_116_116 = in_A[116] & in_B[116];
  assign nP_116_116 = in_A[116] ^ in_B[116];
  assign nG_117_117 = in_A[117] & in_B[117];
  assign nP_117_117 = in_A[117] ^ in_B[117];
  assign nG_118_118 = in_A[118] & in_B[118];
  assign nP_118_118 = in_A[118] ^ in_B[118];
  assign nG_119_119 = in_A[119] & in_B[119];
  assign nP_119_119 = in_A[119] ^ in_B[119];
  assign nG_120_120 = in_A[120] & in_B[120];
  assign nP_120_120 = in_A[120] ^ in_B[120];
  assign nG_121_121 = in_A[121] & in_B[121];
  assign nP_121_121 = in_A[121] ^ in_B[121];
  assign nG_122_122 = in_A[122] & in_B[122];
  assign nP_122_122 = in_A[122] ^ in_B[122];
  assign nG_123_123 = in_A[123] & in_B[123];
  assign nP_123_123 = in_A[123] ^ in_B[123];
  assign nG_124_124 = in_A[124] & in_B[124];
  assign nP_124_124 = in_A[124] ^ in_B[124];
  assign nG_125_125 = in_A[125] & in_B[125];
  assign nP_125_125 = in_A[125] ^ in_B[125];
  assign nG_126_126 = in_A[126] & in_B[126];
  assign nP_126_126 = in_A[126] ^ in_B[126];
  assign nG_127_127 = in_A[127] & in_B[127];
  assign nP_127_127 = in_A[127] ^ in_B[127];
  assign nG_128_128 = in_A[128] & in_B[128];
  assign nP_128_128 = in_A[128] ^ in_B[128];
  assign nG_129_129 = in_A[129] & in_B[129];
  assign nP_129_129 = in_A[129] ^ in_B[129];
  assign nG_130_130 = in_A[130] & in_B[130];
  assign nP_130_130 = in_A[130] ^ in_B[130];
  assign nG_131_131 = in_A[131] & in_B[131];
  assign nP_131_131 = in_A[131] ^ in_B[131];
  assign nG_132_132 = in_A[132] & in_B[132];
  assign nP_132_132 = in_A[132] ^ in_B[132];
  assign nG_133_133 = in_A[133] & in_B[133];
  assign nP_133_133 = in_A[133] ^ in_B[133];
  assign nG_134_134 = in_A[134] & in_B[134];
  assign nP_134_134 = in_A[134] ^ in_B[134];
  assign nG_135_135 = in_A[135] & in_B[135];
  assign nP_135_135 = in_A[135] ^ in_B[135];
  assign nG_136_136 = in_A[136] & in_B[136];
  assign nP_136_136 = in_A[136] ^ in_B[136];
  assign nG_137_137 = in_A[137] & in_B[137];
  assign nP_137_137 = in_A[137] ^ in_B[137];
  assign nG_138_138 = in_A[138] & in_B[138];
  assign nP_138_138 = in_A[138] ^ in_B[138];
  assign nG_139_139 = in_A[139] & in_B[139];
  assign nP_139_139 = in_A[139] ^ in_B[139];
  assign nG_140_140 = in_A[140] & in_B[140];
  assign nP_140_140 = in_A[140] ^ in_B[140];
  assign nG_141_141 = in_A[141] & in_B[141];
  assign nP_141_141 = in_A[141] ^ in_B[141];
  assign nG_142_142 = in_A[142] & in_B[142];
  assign nP_142_142 = in_A[142] ^ in_B[142];
  assign nG_143_143 = in_A[143] & in_B[143];
  assign nP_143_143 = in_A[143] ^ in_B[143];
  assign nG_144_144 = in_A[144] & in_B[144];
  assign nP_144_144 = in_A[144] ^ in_B[144];
  assign nG_145_145 = in_A[145] & in_B[145];
  assign nP_145_145 = in_A[145] ^ in_B[145];
  assign nG_146_146 = in_A[146] & in_B[146];
  assign nP_146_146 = in_A[146] ^ in_B[146];
  assign nG_147_147 = in_A[147] & in_B[147];
  assign nP_147_147 = in_A[147] ^ in_B[147];
  assign nG_148_148 = in_A[148] & in_B[148];
  assign nP_148_148 = in_A[148] ^ in_B[148];
  assign nG_149_149 = in_A[149] & in_B[149];
  assign nP_149_149 = in_A[149] ^ in_B[149];
  assign nG_150_150 = in_A[150] & in_B[150];
  assign nP_150_150 = in_A[150] ^ in_B[150];
  assign nG_151_151 = in_A[151] & in_B[151];
  assign nP_151_151 = in_A[151] ^ in_B[151];
  assign nG_152_152 = in_A[152] & in_B[152];
  assign nP_152_152 = in_A[152] ^ in_B[152];
  assign nG_153_153 = in_A[153] & in_B[153];
  assign nP_153_153 = in_A[153] ^ in_B[153];
  assign nG_154_154 = in_A[154] & in_B[154];
  assign nP_154_154 = in_A[154] ^ in_B[154];
  assign nG_155_155 = in_A[155] & in_B[155];
  assign nP_155_155 = in_A[155] ^ in_B[155];
  assign nG_156_156 = in_A[156] & in_B[156];
  assign nP_156_156 = in_A[156] ^ in_B[156];
  assign nG_157_157 = in_A[157] & in_B[157];
  assign nP_157_157 = in_A[157] ^ in_B[157];
  assign nG_158_158 = in_A[158] & in_B[158];
  assign nP_158_158 = in_A[158] ^ in_B[158];
  assign nG_159_159 = in_A[159] & in_B[159];
  assign nP_159_159 = in_A[159] ^ in_B[159];
  assign nG_160_160 = in_A[160] & in_B[160];
  assign nP_160_160 = in_A[160] ^ in_B[160];
  assign nG_161_161 = in_A[161] & in_B[161];
  assign nP_161_161 = in_A[161] ^ in_B[161];
  assign nG_162_162 = in_A[162] & in_B[162];
  assign nP_162_162 = in_A[162] ^ in_B[162];
  assign nG_163_163 = in_A[163] & in_B[163];
  assign nP_163_163 = in_A[163] ^ in_B[163];
  assign nG_164_164 = in_A[164] & in_B[164];
  assign nP_164_164 = in_A[164] ^ in_B[164];
  assign nG_165_165 = in_A[165] & in_B[165];
  assign nP_165_165 = in_A[165] ^ in_B[165];
  assign nG_166_166 = in_A[166] & in_B[166];
  assign nP_166_166 = in_A[166] ^ in_B[166];
  assign nG_167_167 = in_A[167] & in_B[167];
  assign nP_167_167 = in_A[167] ^ in_B[167];
  assign nG_168_168 = in_A[168] & in_B[168];
  assign nP_168_168 = in_A[168] ^ in_B[168];
  assign nG_169_169 = in_A[169] & in_B[169];
  assign nP_169_169 = in_A[169] ^ in_B[169];
  assign nG_170_170 = in_A[170] & in_B[170];
  assign nP_170_170 = in_A[170] ^ in_B[170];
  assign nG_171_171 = in_A[171] & in_B[171];
  assign nP_171_171 = in_A[171] ^ in_B[171];
  assign nG_172_172 = in_A[172] & in_B[172];
  assign nP_172_172 = in_A[172] ^ in_B[172];
  assign nG_173_173 = in_A[173] & in_B[173];
  assign nP_173_173 = in_A[173] ^ in_B[173];
  assign nG_174_174 = in_A[174] & in_B[174];
  assign nP_174_174 = in_A[174] ^ in_B[174];
  assign nG_175_175 = in_A[175] & in_B[175];
  assign nP_175_175 = in_A[175] ^ in_B[175];
  assign nG_176_176 = in_A[176] & in_B[176];
  assign nP_176_176 = in_A[176] ^ in_B[176];
  assign nG_177_177 = in_A[177] & in_B[177];
  assign nP_177_177 = in_A[177] ^ in_B[177];
  assign nG_178_178 = in_A[178] & in_B[178];
  assign nP_178_178 = in_A[178] ^ in_B[178];
  assign nG_179_179 = in_A[179] & in_B[179];
  assign nP_179_179 = in_A[179] ^ in_B[179];
  assign nG_180_180 = in_A[180] & in_B[180];
  assign nP_180_180 = in_A[180] ^ in_B[180];
  assign nG_181_181 = in_A[181] & in_B[181];
  assign nP_181_181 = in_A[181] ^ in_B[181];
  assign nG_182_182 = in_A[182] & in_B[182];
  assign nP_182_182 = in_A[182] ^ in_B[182];
  assign nG_183_183 = in_A[183] & in_B[183];
  assign nP_183_183 = in_A[183] ^ in_B[183];
  assign nG_184_184 = in_A[184] & in_B[184];
  assign nP_184_184 = in_A[184] ^ in_B[184];
  assign nG_185_185 = in_A[185] & in_B[185];
  assign nP_185_185 = in_A[185] ^ in_B[185];
  assign nG_186_186 = in_A[186] & in_B[186];
  assign nP_186_186 = in_A[186] ^ in_B[186];
  assign nG_187_187 = in_A[187] & in_B[187];
  assign nP_187_187 = in_A[187] ^ in_B[187];
  assign nG_188_188 = in_A[188] & in_B[188];
  assign nP_188_188 = in_A[188] ^ in_B[188];
  assign nG_189_189 = in_A[189] & in_B[189];
  assign nP_189_189 = in_A[189] ^ in_B[189];
  assign nG_190_190 = in_A[190] & in_B[190];
  assign nP_190_190 = in_A[190] ^ in_B[190];
  assign nG_191_191 = in_A[191] & in_B[191];
  assign nP_191_191 = in_A[191] ^ in_B[191];
  assign nG_192_192 = in_A[192] & in_B[192];
  assign nP_192_192 = in_A[192] ^ in_B[192];
  assign nG_193_193 = in_A[193] & in_B[193];
  assign nP_193_193 = in_A[193] ^ in_B[193];
  assign nG_194_194 = in_A[194] & in_B[194];
  assign nP_194_194 = in_A[194] ^ in_B[194];
  assign nG_195_195 = in_A[195] & in_B[195];
  assign nP_195_195 = in_A[195] ^ in_B[195];
  assign nG_196_196 = in_A[196] & in_B[196];
  assign nP_196_196 = in_A[196] ^ in_B[196];
  assign nG_197_197 = in_A[197] & in_B[197];
  assign nP_197_197 = in_A[197] ^ in_B[197];
  assign nG_198_198 = in_A[198] & in_B[198];
  assign nP_198_198 = in_A[198] ^ in_B[198];
  assign nG_199_199 = in_A[199] & in_B[199];
  assign nP_199_199 = in_A[199] ^ in_B[199];
  assign nG_200_200 = in_A[200] & in_B[200];
  assign nP_200_200 = in_A[200] ^ in_B[200];
  assign nG_201_201 = in_A[201] & in_B[201];
  assign nP_201_201 = in_A[201] ^ in_B[201];
  assign nG_202_202 = in_A[202] & in_B[202];
  assign nP_202_202 = in_A[202] ^ in_B[202];
  assign nG_203_203 = in_A[203] & in_B[203];
  assign nP_203_203 = in_A[203] ^ in_B[203];
  assign nG_204_204 = in_A[204] & in_B[204];
  assign nP_204_204 = in_A[204] ^ in_B[204];
  assign nG_205_205 = in_A[205] & in_B[205];
  assign nP_205_205 = in_A[205] ^ in_B[205];
  assign nG_206_206 = in_A[206] & in_B[206];
  assign nP_206_206 = in_A[206] ^ in_B[206];
  assign nG_207_207 = in_A[207] & in_B[207];
  assign nP_207_207 = in_A[207] ^ in_B[207];
  assign nG_208_208 = in_A[208] & in_B[208];
  assign nP_208_208 = in_A[208] ^ in_B[208];
  assign nG_209_209 = in_A[209] & in_B[209];
  assign nP_209_209 = in_A[209] ^ in_B[209];
  assign nG_210_210 = in_A[210] & in_B[210];
  assign nP_210_210 = in_A[210] ^ in_B[210];
  assign nG_211_211 = in_A[211] & in_B[211];
  assign nP_211_211 = in_A[211] ^ in_B[211];
  assign nG_212_212 = in_A[212] & in_B[212];
  assign nP_212_212 = in_A[212] ^ in_B[212];
  assign nG_213_213 = in_A[213] & in_B[213];
  assign nP_213_213 = in_A[213] ^ in_B[213];
  assign nG_214_214 = in_A[214] & in_B[214];
  assign nP_214_214 = in_A[214] ^ in_B[214];
  assign nG_215_215 = in_A[215] & in_B[215];
  assign nP_215_215 = in_A[215] ^ in_B[215];
  assign nG_216_216 = in_A[216] & in_B[216];
  assign nP_216_216 = in_A[216] ^ in_B[216];
  assign nG_217_217 = in_A[217] & in_B[217];
  assign nP_217_217 = in_A[217] ^ in_B[217];
  assign nG_218_218 = in_A[218] & in_B[218];
  assign nP_218_218 = in_A[218] ^ in_B[218];
  assign nG_219_219 = in_A[219] & in_B[219];
  assign nP_219_219 = in_A[219] ^ in_B[219];
  assign nG_220_220 = in_A[220] & in_B[220];
  assign nP_220_220 = in_A[220] ^ in_B[220];
  assign nG_221_221 = in_A[221] & in_B[221];
  assign nP_221_221 = in_A[221] ^ in_B[221];
  assign nG_222_222 = in_A[222] & in_B[222];
  assign nP_222_222 = in_A[222] ^ in_B[222];
  assign nG_223_223 = in_A[223] & in_B[223];
  assign nP_223_223 = in_A[223] ^ in_B[223];
  assign nG_224_224 = in_A[224] & in_B[224];
  assign nP_224_224 = in_A[224] ^ in_B[224];
  assign nG_225_225 = in_A[225] & in_B[225];
  assign nP_225_225 = in_A[225] ^ in_B[225];
  assign nG_226_226 = in_A[226] & in_B[226];
  assign nP_226_226 = in_A[226] ^ in_B[226];
  assign nG_227_227 = in_A[227] & in_B[227];
  assign nP_227_227 = in_A[227] ^ in_B[227];
  assign nG_228_228 = in_A[228] & in_B[228];
  assign nP_228_228 = in_A[228] ^ in_B[228];
  assign nG_229_229 = in_A[229] & in_B[229];
  assign nP_229_229 = in_A[229] ^ in_B[229];
  assign nG_230_230 = in_A[230] & in_B[230];
  assign nP_230_230 = in_A[230] ^ in_B[230];
  assign nG_231_231 = in_A[231] & in_B[231];
  assign nP_231_231 = in_A[231] ^ in_B[231];
  assign nG_232_232 = in_A[232] & in_B[232];
  assign nP_232_232 = in_A[232] ^ in_B[232];
  assign nG_233_233 = in_A[233] & in_B[233];
  assign nP_233_233 = in_A[233] ^ in_B[233];
  assign nG_234_234 = in_A[234] & in_B[234];
  assign nP_234_234 = in_A[234] ^ in_B[234];
  assign nG_235_235 = in_A[235] & in_B[235];
  assign nP_235_235 = in_A[235] ^ in_B[235];
  assign nG_236_236 = in_A[236] & in_B[236];
  assign nP_236_236 = in_A[236] ^ in_B[236];
  assign nG_237_237 = in_A[237] & in_B[237];
  assign nP_237_237 = in_A[237] ^ in_B[237];
  assign nG_238_238 = in_A[238] & in_B[238];
  assign nP_238_238 = in_A[238] ^ in_B[238];
  assign nG_239_239 = in_A[239] & in_B[239];
  assign nP_239_239 = in_A[239] ^ in_B[239];
  assign nG_240_240 = in_A[240] & in_B[240];
  assign nP_240_240 = in_A[240] ^ in_B[240];
  assign nG_241_241 = in_A[241] & in_B[241];
  assign nP_241_241 = in_A[241] ^ in_B[241];
  assign nG_242_242 = in_A[242] & in_B[242];
  assign nP_242_242 = in_A[242] ^ in_B[242];
  assign nG_243_243 = in_A[243] & in_B[243];
  assign nP_243_243 = in_A[243] ^ in_B[243];
  assign nG_244_244 = in_A[244] & in_B[244];
  assign nP_244_244 = in_A[244] ^ in_B[244];
  assign nG_245_245 = in_A[245] & in_B[245];
  assign nP_245_245 = in_A[245] ^ in_B[245];
  assign nG_246_246 = in_A[246] & in_B[246];
  assign nP_246_246 = in_A[246] ^ in_B[246];
  assign nG_247_247 = in_A[247] & in_B[247];
  assign nP_247_247 = in_A[247] ^ in_B[247];
  assign nG_248_248 = in_A[248] & in_B[248];
  assign nP_248_248 = in_A[248] ^ in_B[248];
  assign nG_249_249 = in_A[249] & in_B[249];
  assign nP_249_249 = in_A[249] ^ in_B[249];
  assign nG_250_250 = in_A[250] & in_B[250];
  assign nP_250_250 = in_A[250] ^ in_B[250];
  assign nG_251_251 = in_A[251] & in_B[251];
  assign nP_251_251 = in_A[251] ^ in_B[251];
  assign nG_252_252 = in_A[252] & in_B[252];
  assign nP_252_252 = in_A[252] ^ in_B[252];
  assign nG_253_253 = in_A[253] & in_B[253];
  assign nP_253_253 = in_A[253] ^ in_B[253];
  assign nG_254_254 = in_A[254] & in_B[254];
  assign nP_254_254 = in_A[254] ^ in_B[254];
  assign nG_255_255 = in_A[255] & in_B[255];
  assign nP_255_255 = in_A[255] ^ in_B[255];

  assign nG_255_254 = nG_255_255 | (nP_255_255 & nG_254_254);
  assign nP_255_254 = nP_255_255 & nP_254_254;
  assign nG_254_253 = nG_254_254 | (nP_254_254 & nG_253_253);
  assign nP_254_253 = nP_254_254 & nP_253_253;
  assign nG_253_252 = nG_253_253 | (nP_253_253 & nG_252_252);
  assign nP_253_252 = nP_253_253 & nP_252_252;
  assign nG_252_251 = nG_252_252 | (nP_252_252 & nG_251_251);
  assign nP_252_251 = nP_252_252 & nP_251_251;
  assign nG_251_250 = nG_251_251 | (nP_251_251 & nG_250_250);
  assign nP_251_250 = nP_251_251 & nP_250_250;
  assign nG_250_249 = nG_250_250 | (nP_250_250 & nG_249_249);
  assign nP_250_249 = nP_250_250 & nP_249_249;
  assign nG_249_248 = nG_249_249 | (nP_249_249 & nG_248_248);
  assign nP_249_248 = nP_249_249 & nP_248_248;
  assign nG_248_247 = nG_248_248 | (nP_248_248 & nG_247_247);
  assign nP_248_247 = nP_248_248 & nP_247_247;
  assign nG_247_246 = nG_247_247 | (nP_247_247 & nG_246_246);
  assign nP_247_246 = nP_247_247 & nP_246_246;
  assign nG_246_245 = nG_246_246 | (nP_246_246 & nG_245_245);
  assign nP_246_245 = nP_246_246 & nP_245_245;
  assign nG_245_244 = nG_245_245 | (nP_245_245 & nG_244_244);
  assign nP_245_244 = nP_245_245 & nP_244_244;
  assign nG_244_243 = nG_244_244 | (nP_244_244 & nG_243_243);
  assign nP_244_243 = nP_244_244 & nP_243_243;
  assign nG_243_242 = nG_243_243 | (nP_243_243 & nG_242_242);
  assign nP_243_242 = nP_243_243 & nP_242_242;
  assign nG_242_241 = nG_242_242 | (nP_242_242 & nG_241_241);
  assign nP_242_241 = nP_242_242 & nP_241_241;
  assign nG_241_240 = nG_241_241 | (nP_241_241 & nG_240_240);
  assign nP_241_240 = nP_241_241 & nP_240_240;
  assign nG_240_239 = nG_240_240 | (nP_240_240 & nG_239_239);
  assign nP_240_239 = nP_240_240 & nP_239_239;
  assign nG_239_238 = nG_239_239 | (nP_239_239 & nG_238_238);
  assign nP_239_238 = nP_239_239 & nP_238_238;
  assign nG_238_237 = nG_238_238 | (nP_238_238 & nG_237_237);
  assign nP_238_237 = nP_238_238 & nP_237_237;
  assign nG_237_236 = nG_237_237 | (nP_237_237 & nG_236_236);
  assign nP_237_236 = nP_237_237 & nP_236_236;
  assign nG_236_235 = nG_236_236 | (nP_236_236 & nG_235_235);
  assign nP_236_235 = nP_236_236 & nP_235_235;
  assign nG_235_234 = nG_235_235 | (nP_235_235 & nG_234_234);
  assign nP_235_234 = nP_235_235 & nP_234_234;
  assign nG_234_233 = nG_234_234 | (nP_234_234 & nG_233_233);
  assign nP_234_233 = nP_234_234 & nP_233_233;
  assign nG_233_232 = nG_233_233 | (nP_233_233 & nG_232_232);
  assign nP_233_232 = nP_233_233 & nP_232_232;
  assign nG_232_231 = nG_232_232 | (nP_232_232 & nG_231_231);
  assign nP_232_231 = nP_232_232 & nP_231_231;
  assign nG_231_230 = nG_231_231 | (nP_231_231 & nG_230_230);
  assign nP_231_230 = nP_231_231 & nP_230_230;
  assign nG_230_229 = nG_230_230 | (nP_230_230 & nG_229_229);
  assign nP_230_229 = nP_230_230 & nP_229_229;
  assign nG_229_228 = nG_229_229 | (nP_229_229 & nG_228_228);
  assign nP_229_228 = nP_229_229 & nP_228_228;
  assign nG_228_227 = nG_228_228 | (nP_228_228 & nG_227_227);
  assign nP_228_227 = nP_228_228 & nP_227_227;
  assign nG_227_226 = nG_227_227 | (nP_227_227 & nG_226_226);
  assign nP_227_226 = nP_227_227 & nP_226_226;
  assign nG_226_225 = nG_226_226 | (nP_226_226 & nG_225_225);
  assign nP_226_225 = nP_226_226 & nP_225_225;
  assign nG_225_224 = nG_225_225 | (nP_225_225 & nG_224_224);
  assign nP_225_224 = nP_225_225 & nP_224_224;
  assign nG_224_223 = nG_224_224 | (nP_224_224 & nG_223_223);
  assign nP_224_223 = nP_224_224 & nP_223_223;
  assign nG_223_222 = nG_223_223 | (nP_223_223 & nG_222_222);
  assign nP_223_222 = nP_223_223 & nP_222_222;
  assign nG_222_221 = nG_222_222 | (nP_222_222 & nG_221_221);
  assign nP_222_221 = nP_222_222 & nP_221_221;
  assign nG_221_220 = nG_221_221 | (nP_221_221 & nG_220_220);
  assign nP_221_220 = nP_221_221 & nP_220_220;
  assign nG_220_219 = nG_220_220 | (nP_220_220 & nG_219_219);
  assign nP_220_219 = nP_220_220 & nP_219_219;
  assign nG_219_218 = nG_219_219 | (nP_219_219 & nG_218_218);
  assign nP_219_218 = nP_219_219 & nP_218_218;
  assign nG_218_217 = nG_218_218 | (nP_218_218 & nG_217_217);
  assign nP_218_217 = nP_218_218 & nP_217_217;
  assign nG_217_216 = nG_217_217 | (nP_217_217 & nG_216_216);
  assign nP_217_216 = nP_217_217 & nP_216_216;
  assign nG_216_215 = nG_216_216 | (nP_216_216 & nG_215_215);
  assign nP_216_215 = nP_216_216 & nP_215_215;
  assign nG_215_214 = nG_215_215 | (nP_215_215 & nG_214_214);
  assign nP_215_214 = nP_215_215 & nP_214_214;
  assign nG_214_213 = nG_214_214 | (nP_214_214 & nG_213_213);
  assign nP_214_213 = nP_214_214 & nP_213_213;
  assign nG_213_212 = nG_213_213 | (nP_213_213 & nG_212_212);
  assign nP_213_212 = nP_213_213 & nP_212_212;
  assign nG_212_211 = nG_212_212 | (nP_212_212 & nG_211_211);
  assign nP_212_211 = nP_212_212 & nP_211_211;
  assign nG_211_210 = nG_211_211 | (nP_211_211 & nG_210_210);
  assign nP_211_210 = nP_211_211 & nP_210_210;
  assign nG_210_209 = nG_210_210 | (nP_210_210 & nG_209_209);
  assign nP_210_209 = nP_210_210 & nP_209_209;
  assign nG_209_208 = nG_209_209 | (nP_209_209 & nG_208_208);
  assign nP_209_208 = nP_209_209 & nP_208_208;
  assign nG_208_207 = nG_208_208 | (nP_208_208 & nG_207_207);
  assign nP_208_207 = nP_208_208 & nP_207_207;
  assign nG_207_206 = nG_207_207 | (nP_207_207 & nG_206_206);
  assign nP_207_206 = nP_207_207 & nP_206_206;
  assign nG_206_205 = nG_206_206 | (nP_206_206 & nG_205_205);
  assign nP_206_205 = nP_206_206 & nP_205_205;
  assign nG_205_204 = nG_205_205 | (nP_205_205 & nG_204_204);
  assign nP_205_204 = nP_205_205 & nP_204_204;
  assign nG_204_203 = nG_204_204 | (nP_204_204 & nG_203_203);
  assign nP_204_203 = nP_204_204 & nP_203_203;
  assign nG_203_202 = nG_203_203 | (nP_203_203 & nG_202_202);
  assign nP_203_202 = nP_203_203 & nP_202_202;
  assign nG_202_201 = nG_202_202 | (nP_202_202 & nG_201_201);
  assign nP_202_201 = nP_202_202 & nP_201_201;
  assign nG_201_200 = nG_201_201 | (nP_201_201 & nG_200_200);
  assign nP_201_200 = nP_201_201 & nP_200_200;
  assign nG_200_199 = nG_200_200 | (nP_200_200 & nG_199_199);
  assign nP_200_199 = nP_200_200 & nP_199_199;
  assign nG_199_198 = nG_199_199 | (nP_199_199 & nG_198_198);
  assign nP_199_198 = nP_199_199 & nP_198_198;
  assign nG_198_197 = nG_198_198 | (nP_198_198 & nG_197_197);
  assign nP_198_197 = nP_198_198 & nP_197_197;
  assign nG_197_196 = nG_197_197 | (nP_197_197 & nG_196_196);
  assign nP_197_196 = nP_197_197 & nP_196_196;
  assign nG_196_195 = nG_196_196 | (nP_196_196 & nG_195_195);
  assign nP_196_195 = nP_196_196 & nP_195_195;
  assign nG_195_194 = nG_195_195 | (nP_195_195 & nG_194_194);
  assign nP_195_194 = nP_195_195 & nP_194_194;
  assign nG_194_193 = nG_194_194 | (nP_194_194 & nG_193_193);
  assign nP_194_193 = nP_194_194 & nP_193_193;
  assign nG_193_192 = nG_193_193 | (nP_193_193 & nG_192_192);
  assign nP_193_192 = nP_193_193 & nP_192_192;
  assign nG_192_191 = nG_192_192 | (nP_192_192 & nG_191_191);
  assign nP_192_191 = nP_192_192 & nP_191_191;
  assign nG_191_190 = nG_191_191 | (nP_191_191 & nG_190_190);
  assign nP_191_190 = nP_191_191 & nP_190_190;
  assign nG_190_189 = nG_190_190 | (nP_190_190 & nG_189_189);
  assign nP_190_189 = nP_190_190 & nP_189_189;
  assign nG_189_188 = nG_189_189 | (nP_189_189 & nG_188_188);
  assign nP_189_188 = nP_189_189 & nP_188_188;
  assign nG_188_187 = nG_188_188 | (nP_188_188 & nG_187_187);
  assign nP_188_187 = nP_188_188 & nP_187_187;
  assign nG_187_186 = nG_187_187 | (nP_187_187 & nG_186_186);
  assign nP_187_186 = nP_187_187 & nP_186_186;
  assign nG_186_185 = nG_186_186 | (nP_186_186 & nG_185_185);
  assign nP_186_185 = nP_186_186 & nP_185_185;
  assign nG_185_184 = nG_185_185 | (nP_185_185 & nG_184_184);
  assign nP_185_184 = nP_185_185 & nP_184_184;
  assign nG_184_183 = nG_184_184 | (nP_184_184 & nG_183_183);
  assign nP_184_183 = nP_184_184 & nP_183_183;
  assign nG_183_182 = nG_183_183 | (nP_183_183 & nG_182_182);
  assign nP_183_182 = nP_183_183 & nP_182_182;
  assign nG_182_181 = nG_182_182 | (nP_182_182 & nG_181_181);
  assign nP_182_181 = nP_182_182 & nP_181_181;
  assign nG_181_180 = nG_181_181 | (nP_181_181 & nG_180_180);
  assign nP_181_180 = nP_181_181 & nP_180_180;
  assign nG_180_179 = nG_180_180 | (nP_180_180 & nG_179_179);
  assign nP_180_179 = nP_180_180 & nP_179_179;
  assign nG_179_178 = nG_179_179 | (nP_179_179 & nG_178_178);
  assign nP_179_178 = nP_179_179 & nP_178_178;
  assign nG_178_177 = nG_178_178 | (nP_178_178 & nG_177_177);
  assign nP_178_177 = nP_178_178 & nP_177_177;
  assign nG_177_176 = nG_177_177 | (nP_177_177 & nG_176_176);
  assign nP_177_176 = nP_177_177 & nP_176_176;
  assign nG_176_175 = nG_176_176 | (nP_176_176 & nG_175_175);
  assign nP_176_175 = nP_176_176 & nP_175_175;
  assign nG_175_174 = nG_175_175 | (nP_175_175 & nG_174_174);
  assign nP_175_174 = nP_175_175 & nP_174_174;
  assign nG_174_173 = nG_174_174 | (nP_174_174 & nG_173_173);
  assign nP_174_173 = nP_174_174 & nP_173_173;
  assign nG_173_172 = nG_173_173 | (nP_173_173 & nG_172_172);
  assign nP_173_172 = nP_173_173 & nP_172_172;
  assign nG_172_171 = nG_172_172 | (nP_172_172 & nG_171_171);
  assign nP_172_171 = nP_172_172 & nP_171_171;
  assign nG_171_170 = nG_171_171 | (nP_171_171 & nG_170_170);
  assign nP_171_170 = nP_171_171 & nP_170_170;
  assign nG_170_169 = nG_170_170 | (nP_170_170 & nG_169_169);
  assign nP_170_169 = nP_170_170 & nP_169_169;
  assign nG_169_168 = nG_169_169 | (nP_169_169 & nG_168_168);
  assign nP_169_168 = nP_169_169 & nP_168_168;
  assign nG_168_167 = nG_168_168 | (nP_168_168 & nG_167_167);
  assign nP_168_167 = nP_168_168 & nP_167_167;
  assign nG_167_166 = nG_167_167 | (nP_167_167 & nG_166_166);
  assign nP_167_166 = nP_167_167 & nP_166_166;
  assign nG_166_165 = nG_166_166 | (nP_166_166 & nG_165_165);
  assign nP_166_165 = nP_166_166 & nP_165_165;
  assign nG_165_164 = nG_165_165 | (nP_165_165 & nG_164_164);
  assign nP_165_164 = nP_165_165 & nP_164_164;
  assign nG_164_163 = nG_164_164 | (nP_164_164 & nG_163_163);
  assign nP_164_163 = nP_164_164 & nP_163_163;
  assign nG_163_162 = nG_163_163 | (nP_163_163 & nG_162_162);
  assign nP_163_162 = nP_163_163 & nP_162_162;
  assign nG_162_161 = nG_162_162 | (nP_162_162 & nG_161_161);
  assign nP_162_161 = nP_162_162 & nP_161_161;
  assign nG_161_160 = nG_161_161 | (nP_161_161 & nG_160_160);
  assign nP_161_160 = nP_161_161 & nP_160_160;
  assign nG_160_159 = nG_160_160 | (nP_160_160 & nG_159_159);
  assign nP_160_159 = nP_160_160 & nP_159_159;
  assign nG_159_158 = nG_159_159 | (nP_159_159 & nG_158_158);
  assign nP_159_158 = nP_159_159 & nP_158_158;
  assign nG_158_157 = nG_158_158 | (nP_158_158 & nG_157_157);
  assign nP_158_157 = nP_158_158 & nP_157_157;
  assign nG_157_156 = nG_157_157 | (nP_157_157 & nG_156_156);
  assign nP_157_156 = nP_157_157 & nP_156_156;
  assign nG_156_155 = nG_156_156 | (nP_156_156 & nG_155_155);
  assign nP_156_155 = nP_156_156 & nP_155_155;
  assign nG_155_154 = nG_155_155 | (nP_155_155 & nG_154_154);
  assign nP_155_154 = nP_155_155 & nP_154_154;
  assign nG_154_153 = nG_154_154 | (nP_154_154 & nG_153_153);
  assign nP_154_153 = nP_154_154 & nP_153_153;
  assign nG_153_152 = nG_153_153 | (nP_153_153 & nG_152_152);
  assign nP_153_152 = nP_153_153 & nP_152_152;
  assign nG_152_151 = nG_152_152 | (nP_152_152 & nG_151_151);
  assign nP_152_151 = nP_152_152 & nP_151_151;
  assign nG_151_150 = nG_151_151 | (nP_151_151 & nG_150_150);
  assign nP_151_150 = nP_151_151 & nP_150_150;
  assign nG_150_149 = nG_150_150 | (nP_150_150 & nG_149_149);
  assign nP_150_149 = nP_150_150 & nP_149_149;
  assign nG_149_148 = nG_149_149 | (nP_149_149 & nG_148_148);
  assign nP_149_148 = nP_149_149 & nP_148_148;
  assign nG_148_147 = nG_148_148 | (nP_148_148 & nG_147_147);
  assign nP_148_147 = nP_148_148 & nP_147_147;
  assign nG_147_146 = nG_147_147 | (nP_147_147 & nG_146_146);
  assign nP_147_146 = nP_147_147 & nP_146_146;
  assign nG_146_145 = nG_146_146 | (nP_146_146 & nG_145_145);
  assign nP_146_145 = nP_146_146 & nP_145_145;
  assign nG_145_144 = nG_145_145 | (nP_145_145 & nG_144_144);
  assign nP_145_144 = nP_145_145 & nP_144_144;
  assign nG_144_143 = nG_144_144 | (nP_144_144 & nG_143_143);
  assign nP_144_143 = nP_144_144 & nP_143_143;
  assign nG_143_142 = nG_143_143 | (nP_143_143 & nG_142_142);
  assign nP_143_142 = nP_143_143 & nP_142_142;
  assign nG_142_141 = nG_142_142 | (nP_142_142 & nG_141_141);
  assign nP_142_141 = nP_142_142 & nP_141_141;
  assign nG_141_140 = nG_141_141 | (nP_141_141 & nG_140_140);
  assign nP_141_140 = nP_141_141 & nP_140_140;
  assign nG_140_139 = nG_140_140 | (nP_140_140 & nG_139_139);
  assign nP_140_139 = nP_140_140 & nP_139_139;
  assign nG_139_138 = nG_139_139 | (nP_139_139 & nG_138_138);
  assign nP_139_138 = nP_139_139 & nP_138_138;
  assign nG_138_137 = nG_138_138 | (nP_138_138 & nG_137_137);
  assign nP_138_137 = nP_138_138 & nP_137_137;
  assign nG_137_136 = nG_137_137 | (nP_137_137 & nG_136_136);
  assign nP_137_136 = nP_137_137 & nP_136_136;
  assign nG_136_135 = nG_136_136 | (nP_136_136 & nG_135_135);
  assign nP_136_135 = nP_136_136 & nP_135_135;
  assign nG_135_134 = nG_135_135 | (nP_135_135 & nG_134_134);
  assign nP_135_134 = nP_135_135 & nP_134_134;
  assign nG_134_133 = nG_134_134 | (nP_134_134 & nG_133_133);
  assign nP_134_133 = nP_134_134 & nP_133_133;
  assign nG_133_132 = nG_133_133 | (nP_133_133 & nG_132_132);
  assign nP_133_132 = nP_133_133 & nP_132_132;
  assign nG_132_131 = nG_132_132 | (nP_132_132 & nG_131_131);
  assign nP_132_131 = nP_132_132 & nP_131_131;
  assign nG_131_130 = nG_131_131 | (nP_131_131 & nG_130_130);
  assign nP_131_130 = nP_131_131 & nP_130_130;
  assign nG_130_129 = nG_130_130 | (nP_130_130 & nG_129_129);
  assign nP_130_129 = nP_130_130 & nP_129_129;
  assign nG_129_128 = nG_129_129 | (nP_129_129 & nG_128_128);
  assign nP_129_128 = nP_129_129 & nP_128_128;
  assign nG_128_127 = nG_128_128 | (nP_128_128 & nG_127_127);
  assign nP_128_127 = nP_128_128 & nP_127_127;
  assign nG_127_126 = nG_127_127 | (nP_127_127 & nG_126_126);
  assign nP_127_126 = nP_127_127 & nP_126_126;
  assign nG_126_125 = nG_126_126 | (nP_126_126 & nG_125_125);
  assign nP_126_125 = nP_126_126 & nP_125_125;
  assign nG_125_124 = nG_125_125 | (nP_125_125 & nG_124_124);
  assign nP_125_124 = nP_125_125 & nP_124_124;
  assign nG_124_123 = nG_124_124 | (nP_124_124 & nG_123_123);
  assign nP_124_123 = nP_124_124 & nP_123_123;
  assign nG_123_122 = nG_123_123 | (nP_123_123 & nG_122_122);
  assign nP_123_122 = nP_123_123 & nP_122_122;
  assign nG_122_121 = nG_122_122 | (nP_122_122 & nG_121_121);
  assign nP_122_121 = nP_122_122 & nP_121_121;
  assign nG_121_120 = nG_121_121 | (nP_121_121 & nG_120_120);
  assign nP_121_120 = nP_121_121 & nP_120_120;
  assign nG_120_119 = nG_120_120 | (nP_120_120 & nG_119_119);
  assign nP_120_119 = nP_120_120 & nP_119_119;
  assign nG_119_118 = nG_119_119 | (nP_119_119 & nG_118_118);
  assign nP_119_118 = nP_119_119 & nP_118_118;
  assign nG_118_117 = nG_118_118 | (nP_118_118 & nG_117_117);
  assign nP_118_117 = nP_118_118 & nP_117_117;
  assign nG_117_116 = nG_117_117 | (nP_117_117 & nG_116_116);
  assign nP_117_116 = nP_117_117 & nP_116_116;
  assign nG_116_115 = nG_116_116 | (nP_116_116 & nG_115_115);
  assign nP_116_115 = nP_116_116 & nP_115_115;
  assign nG_115_114 = nG_115_115 | (nP_115_115 & nG_114_114);
  assign nP_115_114 = nP_115_115 & nP_114_114;
  assign nG_114_113 = nG_114_114 | (nP_114_114 & nG_113_113);
  assign nP_114_113 = nP_114_114 & nP_113_113;
  assign nG_113_112 = nG_113_113 | (nP_113_113 & nG_112_112);
  assign nP_113_112 = nP_113_113 & nP_112_112;
  assign nG_112_111 = nG_112_112 | (nP_112_112 & nG_111_111);
  assign nP_112_111 = nP_112_112 & nP_111_111;
  assign nG_111_110 = nG_111_111 | (nP_111_111 & nG_110_110);
  assign nP_111_110 = nP_111_111 & nP_110_110;
  assign nG_110_109 = nG_110_110 | (nP_110_110 & nG_109_109);
  assign nP_110_109 = nP_110_110 & nP_109_109;
  assign nG_109_108 = nG_109_109 | (nP_109_109 & nG_108_108);
  assign nP_109_108 = nP_109_109 & nP_108_108;
  assign nG_108_107 = nG_108_108 | (nP_108_108 & nG_107_107);
  assign nP_108_107 = nP_108_108 & nP_107_107;
  assign nG_107_106 = nG_107_107 | (nP_107_107 & nG_106_106);
  assign nP_107_106 = nP_107_107 & nP_106_106;
  assign nG_106_105 = nG_106_106 | (nP_106_106 & nG_105_105);
  assign nP_106_105 = nP_106_106 & nP_105_105;
  assign nG_105_104 = nG_105_105 | (nP_105_105 & nG_104_104);
  assign nP_105_104 = nP_105_105 & nP_104_104;
  assign nG_104_103 = nG_104_104 | (nP_104_104 & nG_103_103);
  assign nP_104_103 = nP_104_104 & nP_103_103;
  assign nG_103_102 = nG_103_103 | (nP_103_103 & nG_102_102);
  assign nP_103_102 = nP_103_103 & nP_102_102;
  assign nG_102_101 = nG_102_102 | (nP_102_102 & nG_101_101);
  assign nP_102_101 = nP_102_102 & nP_101_101;
  assign nG_101_100 = nG_101_101 | (nP_101_101 & nG_100_100);
  assign nP_101_100 = nP_101_101 & nP_100_100;
  assign nG_100_99 = nG_100_100 | (nP_100_100 & nG_99_99);
  assign nP_100_99 = nP_100_100 & nP_99_99;
  assign nG_99_98 = nG_99_99 | (nP_99_99 & nG_98_98);
  assign nP_99_98 = nP_99_99 & nP_98_98;
  assign nG_98_97 = nG_98_98 | (nP_98_98 & nG_97_97);
  assign nP_98_97 = nP_98_98 & nP_97_97;
  assign nG_97_96 = nG_97_97 | (nP_97_97 & nG_96_96);
  assign nP_97_96 = nP_97_97 & nP_96_96;
  assign nG_96_95 = nG_96_96 | (nP_96_96 & nG_95_95);
  assign nP_96_95 = nP_96_96 & nP_95_95;
  assign nG_95_94 = nG_95_95 | (nP_95_95 & nG_94_94);
  assign nP_95_94 = nP_95_95 & nP_94_94;
  assign nG_94_93 = nG_94_94 | (nP_94_94 & nG_93_93);
  assign nP_94_93 = nP_94_94 & nP_93_93;
  assign nG_93_92 = nG_93_93 | (nP_93_93 & nG_92_92);
  assign nP_93_92 = nP_93_93 & nP_92_92;
  assign nG_92_91 = nG_92_92 | (nP_92_92 & nG_91_91);
  assign nP_92_91 = nP_92_92 & nP_91_91;
  assign nG_91_90 = nG_91_91 | (nP_91_91 & nG_90_90);
  assign nP_91_90 = nP_91_91 & nP_90_90;
  assign nG_90_89 = nG_90_90 | (nP_90_90 & nG_89_89);
  assign nP_90_89 = nP_90_90 & nP_89_89;
  assign nG_89_88 = nG_89_89 | (nP_89_89 & nG_88_88);
  assign nP_89_88 = nP_89_89 & nP_88_88;
  assign nG_88_87 = nG_88_88 | (nP_88_88 & nG_87_87);
  assign nP_88_87 = nP_88_88 & nP_87_87;
  assign nG_87_86 = nG_87_87 | (nP_87_87 & nG_86_86);
  assign nP_87_86 = nP_87_87 & nP_86_86;
  assign nG_86_85 = nG_86_86 | (nP_86_86 & nG_85_85);
  assign nP_86_85 = nP_86_86 & nP_85_85;
  assign nG_85_84 = nG_85_85 | (nP_85_85 & nG_84_84);
  assign nP_85_84 = nP_85_85 & nP_84_84;
  assign nG_84_83 = nG_84_84 | (nP_84_84 & nG_83_83);
  assign nP_84_83 = nP_84_84 & nP_83_83;
  assign nG_83_82 = nG_83_83 | (nP_83_83 & nG_82_82);
  assign nP_83_82 = nP_83_83 & nP_82_82;
  assign nG_82_81 = nG_82_82 | (nP_82_82 & nG_81_81);
  assign nP_82_81 = nP_82_82 & nP_81_81;
  assign nG_81_80 = nG_81_81 | (nP_81_81 & nG_80_80);
  assign nP_81_80 = nP_81_81 & nP_80_80;
  assign nG_80_79 = nG_80_80 | (nP_80_80 & nG_79_79);
  assign nP_80_79 = nP_80_80 & nP_79_79;
  assign nG_79_78 = nG_79_79 | (nP_79_79 & nG_78_78);
  assign nP_79_78 = nP_79_79 & nP_78_78;
  assign nG_78_77 = nG_78_78 | (nP_78_78 & nG_77_77);
  assign nP_78_77 = nP_78_78 & nP_77_77;
  assign nG_77_76 = nG_77_77 | (nP_77_77 & nG_76_76);
  assign nP_77_76 = nP_77_77 & nP_76_76;
  assign nG_76_75 = nG_76_76 | (nP_76_76 & nG_75_75);
  assign nP_76_75 = nP_76_76 & nP_75_75;
  assign nG_75_74 = nG_75_75 | (nP_75_75 & nG_74_74);
  assign nP_75_74 = nP_75_75 & nP_74_74;
  assign nG_74_73 = nG_74_74 | (nP_74_74 & nG_73_73);
  assign nP_74_73 = nP_74_74 & nP_73_73;
  assign nG_73_72 = nG_73_73 | (nP_73_73 & nG_72_72);
  assign nP_73_72 = nP_73_73 & nP_72_72;
  assign nG_72_71 = nG_72_72 | (nP_72_72 & nG_71_71);
  assign nP_72_71 = nP_72_72 & nP_71_71;
  assign nG_71_70 = nG_71_71 | (nP_71_71 & nG_70_70);
  assign nP_71_70 = nP_71_71 & nP_70_70;
  assign nG_70_69 = nG_70_70 | (nP_70_70 & nG_69_69);
  assign nP_70_69 = nP_70_70 & nP_69_69;
  assign nG_69_68 = nG_69_69 | (nP_69_69 & nG_68_68);
  assign nP_69_68 = nP_69_69 & nP_68_68;
  assign nG_68_67 = nG_68_68 | (nP_68_68 & nG_67_67);
  assign nP_68_67 = nP_68_68 & nP_67_67;
  assign nG_67_66 = nG_67_67 | (nP_67_67 & nG_66_66);
  assign nP_67_66 = nP_67_67 & nP_66_66;
  assign nG_66_65 = nG_66_66 | (nP_66_66 & nG_65_65);
  assign nP_66_65 = nP_66_66 & nP_65_65;
  assign nG_65_64 = nG_65_65 | (nP_65_65 & nG_64_64);
  assign nP_65_64 = nP_65_65 & nP_64_64;
  assign nG_64_63 = nG_64_64 | (nP_64_64 & nG_63_63);
  assign nP_64_63 = nP_64_64 & nP_63_63;
  assign nG_63_62 = nG_63_63 | (nP_63_63 & nG_62_62);
  assign nP_63_62 = nP_63_63 & nP_62_62;
  assign nG_62_61 = nG_62_62 | (nP_62_62 & nG_61_61);
  assign nP_62_61 = nP_62_62 & nP_61_61;
  assign nG_61_60 = nG_61_61 | (nP_61_61 & nG_60_60);
  assign nP_61_60 = nP_61_61 & nP_60_60;
  assign nG_60_59 = nG_60_60 | (nP_60_60 & nG_59_59);
  assign nP_60_59 = nP_60_60 & nP_59_59;
  assign nG_59_58 = nG_59_59 | (nP_59_59 & nG_58_58);
  assign nP_59_58 = nP_59_59 & nP_58_58;
  assign nG_58_57 = nG_58_58 | (nP_58_58 & nG_57_57);
  assign nP_58_57 = nP_58_58 & nP_57_57;
  assign nG_57_56 = nG_57_57 | (nP_57_57 & nG_56_56);
  assign nP_57_56 = nP_57_57 & nP_56_56;
  assign nG_56_55 = nG_56_56 | (nP_56_56 & nG_55_55);
  assign nP_56_55 = nP_56_56 & nP_55_55;
  assign nG_55_54 = nG_55_55 | (nP_55_55 & nG_54_54);
  assign nP_55_54 = nP_55_55 & nP_54_54;
  assign nG_54_53 = nG_54_54 | (nP_54_54 & nG_53_53);
  assign nP_54_53 = nP_54_54 & nP_53_53;
  assign nG_53_52 = nG_53_53 | (nP_53_53 & nG_52_52);
  assign nP_53_52 = nP_53_53 & nP_52_52;
  assign nG_52_51 = nG_52_52 | (nP_52_52 & nG_51_51);
  assign nP_52_51 = nP_52_52 & nP_51_51;
  assign nG_51_50 = nG_51_51 | (nP_51_51 & nG_50_50);
  assign nP_51_50 = nP_51_51 & nP_50_50;
  assign nG_50_49 = nG_50_50 | (nP_50_50 & nG_49_49);
  assign nP_50_49 = nP_50_50 & nP_49_49;
  assign nG_49_48 = nG_49_49 | (nP_49_49 & nG_48_48);
  assign nP_49_48 = nP_49_49 & nP_48_48;
  assign nG_48_47 = nG_48_48 | (nP_48_48 & nG_47_47);
  assign nP_48_47 = nP_48_48 & nP_47_47;
  assign nG_47_46 = nG_47_47 | (nP_47_47 & nG_46_46);
  assign nP_47_46 = nP_47_47 & nP_46_46;
  assign nG_46_45 = nG_46_46 | (nP_46_46 & nG_45_45);
  assign nP_46_45 = nP_46_46 & nP_45_45;
  assign nG_45_44 = nG_45_45 | (nP_45_45 & nG_44_44);
  assign nP_45_44 = nP_45_45 & nP_44_44;
  assign nG_44_43 = nG_44_44 | (nP_44_44 & nG_43_43);
  assign nP_44_43 = nP_44_44 & nP_43_43;
  assign nG_43_42 = nG_43_43 | (nP_43_43 & nG_42_42);
  assign nP_43_42 = nP_43_43 & nP_42_42;
  assign nG_42_41 = nG_42_42 | (nP_42_42 & nG_41_41);
  assign nP_42_41 = nP_42_42 & nP_41_41;
  assign nG_41_40 = nG_41_41 | (nP_41_41 & nG_40_40);
  assign nP_41_40 = nP_41_41 & nP_40_40;
  assign nG_40_39 = nG_40_40 | (nP_40_40 & nG_39_39);
  assign nP_40_39 = nP_40_40 & nP_39_39;
  assign nG_39_38 = nG_39_39 | (nP_39_39 & nG_38_38);
  assign nP_39_38 = nP_39_39 & nP_38_38;
  assign nG_38_37 = nG_38_38 | (nP_38_38 & nG_37_37);
  assign nP_38_37 = nP_38_38 & nP_37_37;
  assign nG_37_36 = nG_37_37 | (nP_37_37 & nG_36_36);
  assign nP_37_36 = nP_37_37 & nP_36_36;
  assign nG_36_35 = nG_36_36 | (nP_36_36 & nG_35_35);
  assign nP_36_35 = nP_36_36 & nP_35_35;
  assign nG_35_34 = nG_35_35 | (nP_35_35 & nG_34_34);
  assign nP_35_34 = nP_35_35 & nP_34_34;
  assign nG_34_33 = nG_34_34 | (nP_34_34 & nG_33_33);
  assign nP_34_33 = nP_34_34 & nP_33_33;
  assign nG_33_32 = nG_33_33 | (nP_33_33 & nG_32_32);
  assign nP_33_32 = nP_33_33 & nP_32_32;
  assign nG_32_31 = nG_32_32 | (nP_32_32 & nG_31_31);
  assign nP_32_31 = nP_32_32 & nP_31_31;
  assign nG_31_30 = nG_31_31 | (nP_31_31 & nG_30_30);
  assign nP_31_30 = nP_31_31 & nP_30_30;
  assign nG_30_29 = nG_30_30 | (nP_30_30 & nG_29_29);
  assign nP_30_29 = nP_30_30 & nP_29_29;
  assign nG_29_28 = nG_29_29 | (nP_29_29 & nG_28_28);
  assign nP_29_28 = nP_29_29 & nP_28_28;
  assign nG_28_27 = nG_28_28 | (nP_28_28 & nG_27_27);
  assign nP_28_27 = nP_28_28 & nP_27_27;
  assign nG_27_26 = nG_27_27 | (nP_27_27 & nG_26_26);
  assign nP_27_26 = nP_27_27 & nP_26_26;
  assign nG_26_25 = nG_26_26 | (nP_26_26 & nG_25_25);
  assign nP_26_25 = nP_26_26 & nP_25_25;
  assign nG_25_24 = nG_25_25 | (nP_25_25 & nG_24_24);
  assign nP_25_24 = nP_25_25 & nP_24_24;
  assign nG_24_23 = nG_24_24 | (nP_24_24 & nG_23_23);
  assign nP_24_23 = nP_24_24 & nP_23_23;
  assign nG_23_22 = nG_23_23 | (nP_23_23 & nG_22_22);
  assign nP_23_22 = nP_23_23 & nP_22_22;
  assign nG_22_21 = nG_22_22 | (nP_22_22 & nG_21_21);
  assign nP_22_21 = nP_22_22 & nP_21_21;
  assign nG_21_20 = nG_21_21 | (nP_21_21 & nG_20_20);
  assign nP_21_20 = nP_21_21 & nP_20_20;
  assign nG_20_19 = nG_20_20 | (nP_20_20 & nG_19_19);
  assign nP_20_19 = nP_20_20 & nP_19_19;
  assign nG_19_18 = nG_19_19 | (nP_19_19 & nG_18_18);
  assign nP_19_18 = nP_19_19 & nP_18_18;
  assign nG_18_17 = nG_18_18 | (nP_18_18 & nG_17_17);
  assign nP_18_17 = nP_18_18 & nP_17_17;
  assign nG_17_16 = nG_17_17 | (nP_17_17 & nG_16_16);
  assign nP_17_16 = nP_17_17 & nP_16_16;
  assign nG_16_15 = nG_16_16 | (nP_16_16 & nG_15_15);
  assign nP_16_15 = nP_16_16 & nP_15_15;
  assign nG_15_14 = nG_15_15 | (nP_15_15 & nG_14_14);
  assign nP_15_14 = nP_15_15 & nP_14_14;
  assign nG_14_13 = nG_14_14 | (nP_14_14 & nG_13_13);
  assign nP_14_13 = nP_14_14 & nP_13_13;
  assign nG_13_12 = nG_13_13 | (nP_13_13 & nG_12_12);
  assign nP_13_12 = nP_13_13 & nP_12_12;
  assign nG_12_11 = nG_12_12 | (nP_12_12 & nG_11_11);
  assign nP_12_11 = nP_12_12 & nP_11_11;
  assign nG_11_10 = nG_11_11 | (nP_11_11 & nG_10_10);
  assign nP_11_10 = nP_11_11 & nP_10_10;
  assign nG_10_9 = nG_10_10 | (nP_10_10 & nG_9_9);
  assign nP_10_9 = nP_10_10 & nP_9_9;
  assign nG_9_8 = nG_9_9 | (nP_9_9 & nG_8_8);
  assign nP_9_8 = nP_9_9 & nP_8_8;
  assign nG_8_7 = nG_8_8 | (nP_8_8 & nG_7_7);
  assign nP_8_7 = nP_8_8 & nP_7_7;
  assign nG_7_6 = nG_7_7 | (nP_7_7 & nG_6_6);
  assign nP_7_6 = nP_7_7 & nP_6_6;
  assign nG_6_5 = nG_6_6 | (nP_6_6 & nG_5_5);
  assign nP_6_5 = nP_6_6 & nP_5_5;
  assign nG_5_4 = nG_5_5 | (nP_5_5 & nG_4_4);
  assign nP_5_4 = nP_5_5 & nP_4_4;
  assign nG_4_3 = nG_4_4 | (nP_4_4 & nG_3_3);
  assign nP_4_3 = nP_4_4 & nP_3_3;
  assign nG_3_2 = nG_3_3 | (nP_3_3 & nG_2_2);
  assign nP_3_2 = nP_3_3 & nP_2_2;
  assign nG_2_1 = nG_2_2 | (nP_2_2 & nG_1_1);
  assign nP_2_1 = nP_2_2 & nP_1_1;
  assign nG_1_0 = nG_1_1 | (nP_1_1 & nG_0_0);
  assign nP_1_0 = nP_1_1 & nP_0_0;

  assign nG_255_252 = nG_255_254 | (nP_255_254 & nG_253_252);
  assign nP_255_252 = nP_255_254 & nP_253_252;
  assign nG_254_251 = nG_254_253 | (nP_254_253 & nG_252_251);
  assign nP_254_251 = nP_254_253 & nP_252_251;
  assign nG_253_250 = nG_253_252 | (nP_253_252 & nG_251_250);
  assign nP_253_250 = nP_253_252 & nP_251_250;
  assign nG_252_249 = nG_252_251 | (nP_252_251 & nG_250_249);
  assign nP_252_249 = nP_252_251 & nP_250_249;
  assign nG_251_248 = nG_251_250 | (nP_251_250 & nG_249_248);
  assign nP_251_248 = nP_251_250 & nP_249_248;
  assign nG_250_247 = nG_250_249 | (nP_250_249 & nG_248_247);
  assign nP_250_247 = nP_250_249 & nP_248_247;
  assign nG_249_246 = nG_249_248 | (nP_249_248 & nG_247_246);
  assign nP_249_246 = nP_249_248 & nP_247_246;
  assign nG_248_245 = nG_248_247 | (nP_248_247 & nG_246_245);
  assign nP_248_245 = nP_248_247 & nP_246_245;
  assign nG_247_244 = nG_247_246 | (nP_247_246 & nG_245_244);
  assign nP_247_244 = nP_247_246 & nP_245_244;
  assign nG_246_243 = nG_246_245 | (nP_246_245 & nG_244_243);
  assign nP_246_243 = nP_246_245 & nP_244_243;
  assign nG_245_242 = nG_245_244 | (nP_245_244 & nG_243_242);
  assign nP_245_242 = nP_245_244 & nP_243_242;
  assign nG_244_241 = nG_244_243 | (nP_244_243 & nG_242_241);
  assign nP_244_241 = nP_244_243 & nP_242_241;
  assign nG_243_240 = nG_243_242 | (nP_243_242 & nG_241_240);
  assign nP_243_240 = nP_243_242 & nP_241_240;
  assign nG_242_239 = nG_242_241 | (nP_242_241 & nG_240_239);
  assign nP_242_239 = nP_242_241 & nP_240_239;
  assign nG_241_238 = nG_241_240 | (nP_241_240 & nG_239_238);
  assign nP_241_238 = nP_241_240 & nP_239_238;
  assign nG_240_237 = nG_240_239 | (nP_240_239 & nG_238_237);
  assign nP_240_237 = nP_240_239 & nP_238_237;
  assign nG_239_236 = nG_239_238 | (nP_239_238 & nG_237_236);
  assign nP_239_236 = nP_239_238 & nP_237_236;
  assign nG_238_235 = nG_238_237 | (nP_238_237 & nG_236_235);
  assign nP_238_235 = nP_238_237 & nP_236_235;
  assign nG_237_234 = nG_237_236 | (nP_237_236 & nG_235_234);
  assign nP_237_234 = nP_237_236 & nP_235_234;
  assign nG_236_233 = nG_236_235 | (nP_236_235 & nG_234_233);
  assign nP_236_233 = nP_236_235 & nP_234_233;
  assign nG_235_232 = nG_235_234 | (nP_235_234 & nG_233_232);
  assign nP_235_232 = nP_235_234 & nP_233_232;
  assign nG_234_231 = nG_234_233 | (nP_234_233 & nG_232_231);
  assign nP_234_231 = nP_234_233 & nP_232_231;
  assign nG_233_230 = nG_233_232 | (nP_233_232 & nG_231_230);
  assign nP_233_230 = nP_233_232 & nP_231_230;
  assign nG_232_229 = nG_232_231 | (nP_232_231 & nG_230_229);
  assign nP_232_229 = nP_232_231 & nP_230_229;
  assign nG_231_228 = nG_231_230 | (nP_231_230 & nG_229_228);
  assign nP_231_228 = nP_231_230 & nP_229_228;
  assign nG_230_227 = nG_230_229 | (nP_230_229 & nG_228_227);
  assign nP_230_227 = nP_230_229 & nP_228_227;
  assign nG_229_226 = nG_229_228 | (nP_229_228 & nG_227_226);
  assign nP_229_226 = nP_229_228 & nP_227_226;
  assign nG_228_225 = nG_228_227 | (nP_228_227 & nG_226_225);
  assign nP_228_225 = nP_228_227 & nP_226_225;
  assign nG_227_224 = nG_227_226 | (nP_227_226 & nG_225_224);
  assign nP_227_224 = nP_227_226 & nP_225_224;
  assign nG_226_223 = nG_226_225 | (nP_226_225 & nG_224_223);
  assign nP_226_223 = nP_226_225 & nP_224_223;
  assign nG_225_222 = nG_225_224 | (nP_225_224 & nG_223_222);
  assign nP_225_222 = nP_225_224 & nP_223_222;
  assign nG_224_221 = nG_224_223 | (nP_224_223 & nG_222_221);
  assign nP_224_221 = nP_224_223 & nP_222_221;
  assign nG_223_220 = nG_223_222 | (nP_223_222 & nG_221_220);
  assign nP_223_220 = nP_223_222 & nP_221_220;
  assign nG_222_219 = nG_222_221 | (nP_222_221 & nG_220_219);
  assign nP_222_219 = nP_222_221 & nP_220_219;
  assign nG_221_218 = nG_221_220 | (nP_221_220 & nG_219_218);
  assign nP_221_218 = nP_221_220 & nP_219_218;
  assign nG_220_217 = nG_220_219 | (nP_220_219 & nG_218_217);
  assign nP_220_217 = nP_220_219 & nP_218_217;
  assign nG_219_216 = nG_219_218 | (nP_219_218 & nG_217_216);
  assign nP_219_216 = nP_219_218 & nP_217_216;
  assign nG_218_215 = nG_218_217 | (nP_218_217 & nG_216_215);
  assign nP_218_215 = nP_218_217 & nP_216_215;
  assign nG_217_214 = nG_217_216 | (nP_217_216 & nG_215_214);
  assign nP_217_214 = nP_217_216 & nP_215_214;
  assign nG_216_213 = nG_216_215 | (nP_216_215 & nG_214_213);
  assign nP_216_213 = nP_216_215 & nP_214_213;
  assign nG_215_212 = nG_215_214 | (nP_215_214 & nG_213_212);
  assign nP_215_212 = nP_215_214 & nP_213_212;
  assign nG_214_211 = nG_214_213 | (nP_214_213 & nG_212_211);
  assign nP_214_211 = nP_214_213 & nP_212_211;
  assign nG_213_210 = nG_213_212 | (nP_213_212 & nG_211_210);
  assign nP_213_210 = nP_213_212 & nP_211_210;
  assign nG_212_209 = nG_212_211 | (nP_212_211 & nG_210_209);
  assign nP_212_209 = nP_212_211 & nP_210_209;
  assign nG_211_208 = nG_211_210 | (nP_211_210 & nG_209_208);
  assign nP_211_208 = nP_211_210 & nP_209_208;
  assign nG_210_207 = nG_210_209 | (nP_210_209 & nG_208_207);
  assign nP_210_207 = nP_210_209 & nP_208_207;
  assign nG_209_206 = nG_209_208 | (nP_209_208 & nG_207_206);
  assign nP_209_206 = nP_209_208 & nP_207_206;
  assign nG_208_205 = nG_208_207 | (nP_208_207 & nG_206_205);
  assign nP_208_205 = nP_208_207 & nP_206_205;
  assign nG_207_204 = nG_207_206 | (nP_207_206 & nG_205_204);
  assign nP_207_204 = nP_207_206 & nP_205_204;
  assign nG_206_203 = nG_206_205 | (nP_206_205 & nG_204_203);
  assign nP_206_203 = nP_206_205 & nP_204_203;
  assign nG_205_202 = nG_205_204 | (nP_205_204 & nG_203_202);
  assign nP_205_202 = nP_205_204 & nP_203_202;
  assign nG_204_201 = nG_204_203 | (nP_204_203 & nG_202_201);
  assign nP_204_201 = nP_204_203 & nP_202_201;
  assign nG_203_200 = nG_203_202 | (nP_203_202 & nG_201_200);
  assign nP_203_200 = nP_203_202 & nP_201_200;
  assign nG_202_199 = nG_202_201 | (nP_202_201 & nG_200_199);
  assign nP_202_199 = nP_202_201 & nP_200_199;
  assign nG_201_198 = nG_201_200 | (nP_201_200 & nG_199_198);
  assign nP_201_198 = nP_201_200 & nP_199_198;
  assign nG_200_197 = nG_200_199 | (nP_200_199 & nG_198_197);
  assign nP_200_197 = nP_200_199 & nP_198_197;
  assign nG_199_196 = nG_199_198 | (nP_199_198 & nG_197_196);
  assign nP_199_196 = nP_199_198 & nP_197_196;
  assign nG_198_195 = nG_198_197 | (nP_198_197 & nG_196_195);
  assign nP_198_195 = nP_198_197 & nP_196_195;
  assign nG_197_194 = nG_197_196 | (nP_197_196 & nG_195_194);
  assign nP_197_194 = nP_197_196 & nP_195_194;
  assign nG_196_193 = nG_196_195 | (nP_196_195 & nG_194_193);
  assign nP_196_193 = nP_196_195 & nP_194_193;
  assign nG_195_192 = nG_195_194 | (nP_195_194 & nG_193_192);
  assign nP_195_192 = nP_195_194 & nP_193_192;
  assign nG_194_191 = nG_194_193 | (nP_194_193 & nG_192_191);
  assign nP_194_191 = nP_194_193 & nP_192_191;
  assign nG_193_190 = nG_193_192 | (nP_193_192 & nG_191_190);
  assign nP_193_190 = nP_193_192 & nP_191_190;
  assign nG_192_189 = nG_192_191 | (nP_192_191 & nG_190_189);
  assign nP_192_189 = nP_192_191 & nP_190_189;
  assign nG_191_188 = nG_191_190 | (nP_191_190 & nG_189_188);
  assign nP_191_188 = nP_191_190 & nP_189_188;
  assign nG_190_187 = nG_190_189 | (nP_190_189 & nG_188_187);
  assign nP_190_187 = nP_190_189 & nP_188_187;
  assign nG_189_186 = nG_189_188 | (nP_189_188 & nG_187_186);
  assign nP_189_186 = nP_189_188 & nP_187_186;
  assign nG_188_185 = nG_188_187 | (nP_188_187 & nG_186_185);
  assign nP_188_185 = nP_188_187 & nP_186_185;
  assign nG_187_184 = nG_187_186 | (nP_187_186 & nG_185_184);
  assign nP_187_184 = nP_187_186 & nP_185_184;
  assign nG_186_183 = nG_186_185 | (nP_186_185 & nG_184_183);
  assign nP_186_183 = nP_186_185 & nP_184_183;
  assign nG_185_182 = nG_185_184 | (nP_185_184 & nG_183_182);
  assign nP_185_182 = nP_185_184 & nP_183_182;
  assign nG_184_181 = nG_184_183 | (nP_184_183 & nG_182_181);
  assign nP_184_181 = nP_184_183 & nP_182_181;
  assign nG_183_180 = nG_183_182 | (nP_183_182 & nG_181_180);
  assign nP_183_180 = nP_183_182 & nP_181_180;
  assign nG_182_179 = nG_182_181 | (nP_182_181 & nG_180_179);
  assign nP_182_179 = nP_182_181 & nP_180_179;
  assign nG_181_178 = nG_181_180 | (nP_181_180 & nG_179_178);
  assign nP_181_178 = nP_181_180 & nP_179_178;
  assign nG_180_177 = nG_180_179 | (nP_180_179 & nG_178_177);
  assign nP_180_177 = nP_180_179 & nP_178_177;
  assign nG_179_176 = nG_179_178 | (nP_179_178 & nG_177_176);
  assign nP_179_176 = nP_179_178 & nP_177_176;
  assign nG_178_175 = nG_178_177 | (nP_178_177 & nG_176_175);
  assign nP_178_175 = nP_178_177 & nP_176_175;
  assign nG_177_174 = nG_177_176 | (nP_177_176 & nG_175_174);
  assign nP_177_174 = nP_177_176 & nP_175_174;
  assign nG_176_173 = nG_176_175 | (nP_176_175 & nG_174_173);
  assign nP_176_173 = nP_176_175 & nP_174_173;
  assign nG_175_172 = nG_175_174 | (nP_175_174 & nG_173_172);
  assign nP_175_172 = nP_175_174 & nP_173_172;
  assign nG_174_171 = nG_174_173 | (nP_174_173 & nG_172_171);
  assign nP_174_171 = nP_174_173 & nP_172_171;
  assign nG_173_170 = nG_173_172 | (nP_173_172 & nG_171_170);
  assign nP_173_170 = nP_173_172 & nP_171_170;
  assign nG_172_169 = nG_172_171 | (nP_172_171 & nG_170_169);
  assign nP_172_169 = nP_172_171 & nP_170_169;
  assign nG_171_168 = nG_171_170 | (nP_171_170 & nG_169_168);
  assign nP_171_168 = nP_171_170 & nP_169_168;
  assign nG_170_167 = nG_170_169 | (nP_170_169 & nG_168_167);
  assign nP_170_167 = nP_170_169 & nP_168_167;
  assign nG_169_166 = nG_169_168 | (nP_169_168 & nG_167_166);
  assign nP_169_166 = nP_169_168 & nP_167_166;
  assign nG_168_165 = nG_168_167 | (nP_168_167 & nG_166_165);
  assign nP_168_165 = nP_168_167 & nP_166_165;
  assign nG_167_164 = nG_167_166 | (nP_167_166 & nG_165_164);
  assign nP_167_164 = nP_167_166 & nP_165_164;
  assign nG_166_163 = nG_166_165 | (nP_166_165 & nG_164_163);
  assign nP_166_163 = nP_166_165 & nP_164_163;
  assign nG_165_162 = nG_165_164 | (nP_165_164 & nG_163_162);
  assign nP_165_162 = nP_165_164 & nP_163_162;
  assign nG_164_161 = nG_164_163 | (nP_164_163 & nG_162_161);
  assign nP_164_161 = nP_164_163 & nP_162_161;
  assign nG_163_160 = nG_163_162 | (nP_163_162 & nG_161_160);
  assign nP_163_160 = nP_163_162 & nP_161_160;
  assign nG_162_159 = nG_162_161 | (nP_162_161 & nG_160_159);
  assign nP_162_159 = nP_162_161 & nP_160_159;
  assign nG_161_158 = nG_161_160 | (nP_161_160 & nG_159_158);
  assign nP_161_158 = nP_161_160 & nP_159_158;
  assign nG_160_157 = nG_160_159 | (nP_160_159 & nG_158_157);
  assign nP_160_157 = nP_160_159 & nP_158_157;
  assign nG_159_156 = nG_159_158 | (nP_159_158 & nG_157_156);
  assign nP_159_156 = nP_159_158 & nP_157_156;
  assign nG_158_155 = nG_158_157 | (nP_158_157 & nG_156_155);
  assign nP_158_155 = nP_158_157 & nP_156_155;
  assign nG_157_154 = nG_157_156 | (nP_157_156 & nG_155_154);
  assign nP_157_154 = nP_157_156 & nP_155_154;
  assign nG_156_153 = nG_156_155 | (nP_156_155 & nG_154_153);
  assign nP_156_153 = nP_156_155 & nP_154_153;
  assign nG_155_152 = nG_155_154 | (nP_155_154 & nG_153_152);
  assign nP_155_152 = nP_155_154 & nP_153_152;
  assign nG_154_151 = nG_154_153 | (nP_154_153 & nG_152_151);
  assign nP_154_151 = nP_154_153 & nP_152_151;
  assign nG_153_150 = nG_153_152 | (nP_153_152 & nG_151_150);
  assign nP_153_150 = nP_153_152 & nP_151_150;
  assign nG_152_149 = nG_152_151 | (nP_152_151 & nG_150_149);
  assign nP_152_149 = nP_152_151 & nP_150_149;
  assign nG_151_148 = nG_151_150 | (nP_151_150 & nG_149_148);
  assign nP_151_148 = nP_151_150 & nP_149_148;
  assign nG_150_147 = nG_150_149 | (nP_150_149 & nG_148_147);
  assign nP_150_147 = nP_150_149 & nP_148_147;
  assign nG_149_146 = nG_149_148 | (nP_149_148 & nG_147_146);
  assign nP_149_146 = nP_149_148 & nP_147_146;
  assign nG_148_145 = nG_148_147 | (nP_148_147 & nG_146_145);
  assign nP_148_145 = nP_148_147 & nP_146_145;
  assign nG_147_144 = nG_147_146 | (nP_147_146 & nG_145_144);
  assign nP_147_144 = nP_147_146 & nP_145_144;
  assign nG_146_143 = nG_146_145 | (nP_146_145 & nG_144_143);
  assign nP_146_143 = nP_146_145 & nP_144_143;
  assign nG_145_142 = nG_145_144 | (nP_145_144 & nG_143_142);
  assign nP_145_142 = nP_145_144 & nP_143_142;
  assign nG_144_141 = nG_144_143 | (nP_144_143 & nG_142_141);
  assign nP_144_141 = nP_144_143 & nP_142_141;
  assign nG_143_140 = nG_143_142 | (nP_143_142 & nG_141_140);
  assign nP_143_140 = nP_143_142 & nP_141_140;
  assign nG_142_139 = nG_142_141 | (nP_142_141 & nG_140_139);
  assign nP_142_139 = nP_142_141 & nP_140_139;
  assign nG_141_138 = nG_141_140 | (nP_141_140 & nG_139_138);
  assign nP_141_138 = nP_141_140 & nP_139_138;
  assign nG_140_137 = nG_140_139 | (nP_140_139 & nG_138_137);
  assign nP_140_137 = nP_140_139 & nP_138_137;
  assign nG_139_136 = nG_139_138 | (nP_139_138 & nG_137_136);
  assign nP_139_136 = nP_139_138 & nP_137_136;
  assign nG_138_135 = nG_138_137 | (nP_138_137 & nG_136_135);
  assign nP_138_135 = nP_138_137 & nP_136_135;
  assign nG_137_134 = nG_137_136 | (nP_137_136 & nG_135_134);
  assign nP_137_134 = nP_137_136 & nP_135_134;
  assign nG_136_133 = nG_136_135 | (nP_136_135 & nG_134_133);
  assign nP_136_133 = nP_136_135 & nP_134_133;
  assign nG_135_132 = nG_135_134 | (nP_135_134 & nG_133_132);
  assign nP_135_132 = nP_135_134 & nP_133_132;
  assign nG_134_131 = nG_134_133 | (nP_134_133 & nG_132_131);
  assign nP_134_131 = nP_134_133 & nP_132_131;
  assign nG_133_130 = nG_133_132 | (nP_133_132 & nG_131_130);
  assign nP_133_130 = nP_133_132 & nP_131_130;
  assign nG_132_129 = nG_132_131 | (nP_132_131 & nG_130_129);
  assign nP_132_129 = nP_132_131 & nP_130_129;
  assign nG_131_128 = nG_131_130 | (nP_131_130 & nG_129_128);
  assign nP_131_128 = nP_131_130 & nP_129_128;
  assign nG_130_127 = nG_130_129 | (nP_130_129 & nG_128_127);
  assign nP_130_127 = nP_130_129 & nP_128_127;
  assign nG_129_126 = nG_129_128 | (nP_129_128 & nG_127_126);
  assign nP_129_126 = nP_129_128 & nP_127_126;
  assign nG_128_125 = nG_128_127 | (nP_128_127 & nG_126_125);
  assign nP_128_125 = nP_128_127 & nP_126_125;
  assign nG_127_124 = nG_127_126 | (nP_127_126 & nG_125_124);
  assign nP_127_124 = nP_127_126 & nP_125_124;
  assign nG_126_123 = nG_126_125 | (nP_126_125 & nG_124_123);
  assign nP_126_123 = nP_126_125 & nP_124_123;
  assign nG_125_122 = nG_125_124 | (nP_125_124 & nG_123_122);
  assign nP_125_122 = nP_125_124 & nP_123_122;
  assign nG_124_121 = nG_124_123 | (nP_124_123 & nG_122_121);
  assign nP_124_121 = nP_124_123 & nP_122_121;
  assign nG_123_120 = nG_123_122 | (nP_123_122 & nG_121_120);
  assign nP_123_120 = nP_123_122 & nP_121_120;
  assign nG_122_119 = nG_122_121 | (nP_122_121 & nG_120_119);
  assign nP_122_119 = nP_122_121 & nP_120_119;
  assign nG_121_118 = nG_121_120 | (nP_121_120 & nG_119_118);
  assign nP_121_118 = nP_121_120 & nP_119_118;
  assign nG_120_117 = nG_120_119 | (nP_120_119 & nG_118_117);
  assign nP_120_117 = nP_120_119 & nP_118_117;
  assign nG_119_116 = nG_119_118 | (nP_119_118 & nG_117_116);
  assign nP_119_116 = nP_119_118 & nP_117_116;
  assign nG_118_115 = nG_118_117 | (nP_118_117 & nG_116_115);
  assign nP_118_115 = nP_118_117 & nP_116_115;
  assign nG_117_114 = nG_117_116 | (nP_117_116 & nG_115_114);
  assign nP_117_114 = nP_117_116 & nP_115_114;
  assign nG_116_113 = nG_116_115 | (nP_116_115 & nG_114_113);
  assign nP_116_113 = nP_116_115 & nP_114_113;
  assign nG_115_112 = nG_115_114 | (nP_115_114 & nG_113_112);
  assign nP_115_112 = nP_115_114 & nP_113_112;
  assign nG_114_111 = nG_114_113 | (nP_114_113 & nG_112_111);
  assign nP_114_111 = nP_114_113 & nP_112_111;
  assign nG_113_110 = nG_113_112 | (nP_113_112 & nG_111_110);
  assign nP_113_110 = nP_113_112 & nP_111_110;
  assign nG_112_109 = nG_112_111 | (nP_112_111 & nG_110_109);
  assign nP_112_109 = nP_112_111 & nP_110_109;
  assign nG_111_108 = nG_111_110 | (nP_111_110 & nG_109_108);
  assign nP_111_108 = nP_111_110 & nP_109_108;
  assign nG_110_107 = nG_110_109 | (nP_110_109 & nG_108_107);
  assign nP_110_107 = nP_110_109 & nP_108_107;
  assign nG_109_106 = nG_109_108 | (nP_109_108 & nG_107_106);
  assign nP_109_106 = nP_109_108 & nP_107_106;
  assign nG_108_105 = nG_108_107 | (nP_108_107 & nG_106_105);
  assign nP_108_105 = nP_108_107 & nP_106_105;
  assign nG_107_104 = nG_107_106 | (nP_107_106 & nG_105_104);
  assign nP_107_104 = nP_107_106 & nP_105_104;
  assign nG_106_103 = nG_106_105 | (nP_106_105 & nG_104_103);
  assign nP_106_103 = nP_106_105 & nP_104_103;
  assign nG_105_102 = nG_105_104 | (nP_105_104 & nG_103_102);
  assign nP_105_102 = nP_105_104 & nP_103_102;
  assign nG_104_101 = nG_104_103 | (nP_104_103 & nG_102_101);
  assign nP_104_101 = nP_104_103 & nP_102_101;
  assign nG_103_100 = nG_103_102 | (nP_103_102 & nG_101_100);
  assign nP_103_100 = nP_103_102 & nP_101_100;
  assign nG_102_99 = nG_102_101 | (nP_102_101 & nG_100_99);
  assign nP_102_99 = nP_102_101 & nP_100_99;
  assign nG_101_98 = nG_101_100 | (nP_101_100 & nG_99_98);
  assign nP_101_98 = nP_101_100 & nP_99_98;
  assign nG_100_97 = nG_100_99 | (nP_100_99 & nG_98_97);
  assign nP_100_97 = nP_100_99 & nP_98_97;
  assign nG_99_96 = nG_99_98 | (nP_99_98 & nG_97_96);
  assign nP_99_96 = nP_99_98 & nP_97_96;
  assign nG_98_95 = nG_98_97 | (nP_98_97 & nG_96_95);
  assign nP_98_95 = nP_98_97 & nP_96_95;
  assign nG_97_94 = nG_97_96 | (nP_97_96 & nG_95_94);
  assign nP_97_94 = nP_97_96 & nP_95_94;
  assign nG_96_93 = nG_96_95 | (nP_96_95 & nG_94_93);
  assign nP_96_93 = nP_96_95 & nP_94_93;
  assign nG_95_92 = nG_95_94 | (nP_95_94 & nG_93_92);
  assign nP_95_92 = nP_95_94 & nP_93_92;
  assign nG_94_91 = nG_94_93 | (nP_94_93 & nG_92_91);
  assign nP_94_91 = nP_94_93 & nP_92_91;
  assign nG_93_90 = nG_93_92 | (nP_93_92 & nG_91_90);
  assign nP_93_90 = nP_93_92 & nP_91_90;
  assign nG_92_89 = nG_92_91 | (nP_92_91 & nG_90_89);
  assign nP_92_89 = nP_92_91 & nP_90_89;
  assign nG_91_88 = nG_91_90 | (nP_91_90 & nG_89_88);
  assign nP_91_88 = nP_91_90 & nP_89_88;
  assign nG_90_87 = nG_90_89 | (nP_90_89 & nG_88_87);
  assign nP_90_87 = nP_90_89 & nP_88_87;
  assign nG_89_86 = nG_89_88 | (nP_89_88 & nG_87_86);
  assign nP_89_86 = nP_89_88 & nP_87_86;
  assign nG_88_85 = nG_88_87 | (nP_88_87 & nG_86_85);
  assign nP_88_85 = nP_88_87 & nP_86_85;
  assign nG_87_84 = nG_87_86 | (nP_87_86 & nG_85_84);
  assign nP_87_84 = nP_87_86 & nP_85_84;
  assign nG_86_83 = nG_86_85 | (nP_86_85 & nG_84_83);
  assign nP_86_83 = nP_86_85 & nP_84_83;
  assign nG_85_82 = nG_85_84 | (nP_85_84 & nG_83_82);
  assign nP_85_82 = nP_85_84 & nP_83_82;
  assign nG_84_81 = nG_84_83 | (nP_84_83 & nG_82_81);
  assign nP_84_81 = nP_84_83 & nP_82_81;
  assign nG_83_80 = nG_83_82 | (nP_83_82 & nG_81_80);
  assign nP_83_80 = nP_83_82 & nP_81_80;
  assign nG_82_79 = nG_82_81 | (nP_82_81 & nG_80_79);
  assign nP_82_79 = nP_82_81 & nP_80_79;
  assign nG_81_78 = nG_81_80 | (nP_81_80 & nG_79_78);
  assign nP_81_78 = nP_81_80 & nP_79_78;
  assign nG_80_77 = nG_80_79 | (nP_80_79 & nG_78_77);
  assign nP_80_77 = nP_80_79 & nP_78_77;
  assign nG_79_76 = nG_79_78 | (nP_79_78 & nG_77_76);
  assign nP_79_76 = nP_79_78 & nP_77_76;
  assign nG_78_75 = nG_78_77 | (nP_78_77 & nG_76_75);
  assign nP_78_75 = nP_78_77 & nP_76_75;
  assign nG_77_74 = nG_77_76 | (nP_77_76 & nG_75_74);
  assign nP_77_74 = nP_77_76 & nP_75_74;
  assign nG_76_73 = nG_76_75 | (nP_76_75 & nG_74_73);
  assign nP_76_73 = nP_76_75 & nP_74_73;
  assign nG_75_72 = nG_75_74 | (nP_75_74 & nG_73_72);
  assign nP_75_72 = nP_75_74 & nP_73_72;
  assign nG_74_71 = nG_74_73 | (nP_74_73 & nG_72_71);
  assign nP_74_71 = nP_74_73 & nP_72_71;
  assign nG_73_70 = nG_73_72 | (nP_73_72 & nG_71_70);
  assign nP_73_70 = nP_73_72 & nP_71_70;
  assign nG_72_69 = nG_72_71 | (nP_72_71 & nG_70_69);
  assign nP_72_69 = nP_72_71 & nP_70_69;
  assign nG_71_68 = nG_71_70 | (nP_71_70 & nG_69_68);
  assign nP_71_68 = nP_71_70 & nP_69_68;
  assign nG_70_67 = nG_70_69 | (nP_70_69 & nG_68_67);
  assign nP_70_67 = nP_70_69 & nP_68_67;
  assign nG_69_66 = nG_69_68 | (nP_69_68 & nG_67_66);
  assign nP_69_66 = nP_69_68 & nP_67_66;
  assign nG_68_65 = nG_68_67 | (nP_68_67 & nG_66_65);
  assign nP_68_65 = nP_68_67 & nP_66_65;
  assign nG_67_64 = nG_67_66 | (nP_67_66 & nG_65_64);
  assign nP_67_64 = nP_67_66 & nP_65_64;
  assign nG_66_63 = nG_66_65 | (nP_66_65 & nG_64_63);
  assign nP_66_63 = nP_66_65 & nP_64_63;
  assign nG_65_62 = nG_65_64 | (nP_65_64 & nG_63_62);
  assign nP_65_62 = nP_65_64 & nP_63_62;
  assign nG_64_61 = nG_64_63 | (nP_64_63 & nG_62_61);
  assign nP_64_61 = nP_64_63 & nP_62_61;
  assign nG_63_60 = nG_63_62 | (nP_63_62 & nG_61_60);
  assign nP_63_60 = nP_63_62 & nP_61_60;
  assign nG_62_59 = nG_62_61 | (nP_62_61 & nG_60_59);
  assign nP_62_59 = nP_62_61 & nP_60_59;
  assign nG_61_58 = nG_61_60 | (nP_61_60 & nG_59_58);
  assign nP_61_58 = nP_61_60 & nP_59_58;
  assign nG_60_57 = nG_60_59 | (nP_60_59 & nG_58_57);
  assign nP_60_57 = nP_60_59 & nP_58_57;
  assign nG_59_56 = nG_59_58 | (nP_59_58 & nG_57_56);
  assign nP_59_56 = nP_59_58 & nP_57_56;
  assign nG_58_55 = nG_58_57 | (nP_58_57 & nG_56_55);
  assign nP_58_55 = nP_58_57 & nP_56_55;
  assign nG_57_54 = nG_57_56 | (nP_57_56 & nG_55_54);
  assign nP_57_54 = nP_57_56 & nP_55_54;
  assign nG_56_53 = nG_56_55 | (nP_56_55 & nG_54_53);
  assign nP_56_53 = nP_56_55 & nP_54_53;
  assign nG_55_52 = nG_55_54 | (nP_55_54 & nG_53_52);
  assign nP_55_52 = nP_55_54 & nP_53_52;
  assign nG_54_51 = nG_54_53 | (nP_54_53 & nG_52_51);
  assign nP_54_51 = nP_54_53 & nP_52_51;
  assign nG_53_50 = nG_53_52 | (nP_53_52 & nG_51_50);
  assign nP_53_50 = nP_53_52 & nP_51_50;
  assign nG_52_49 = nG_52_51 | (nP_52_51 & nG_50_49);
  assign nP_52_49 = nP_52_51 & nP_50_49;
  assign nG_51_48 = nG_51_50 | (nP_51_50 & nG_49_48);
  assign nP_51_48 = nP_51_50 & nP_49_48;
  assign nG_50_47 = nG_50_49 | (nP_50_49 & nG_48_47);
  assign nP_50_47 = nP_50_49 & nP_48_47;
  assign nG_49_46 = nG_49_48 | (nP_49_48 & nG_47_46);
  assign nP_49_46 = nP_49_48 & nP_47_46;
  assign nG_48_45 = nG_48_47 | (nP_48_47 & nG_46_45);
  assign nP_48_45 = nP_48_47 & nP_46_45;
  assign nG_47_44 = nG_47_46 | (nP_47_46 & nG_45_44);
  assign nP_47_44 = nP_47_46 & nP_45_44;
  assign nG_46_43 = nG_46_45 | (nP_46_45 & nG_44_43);
  assign nP_46_43 = nP_46_45 & nP_44_43;
  assign nG_45_42 = nG_45_44 | (nP_45_44 & nG_43_42);
  assign nP_45_42 = nP_45_44 & nP_43_42;
  assign nG_44_41 = nG_44_43 | (nP_44_43 & nG_42_41);
  assign nP_44_41 = nP_44_43 & nP_42_41;
  assign nG_43_40 = nG_43_42 | (nP_43_42 & nG_41_40);
  assign nP_43_40 = nP_43_42 & nP_41_40;
  assign nG_42_39 = nG_42_41 | (nP_42_41 & nG_40_39);
  assign nP_42_39 = nP_42_41 & nP_40_39;
  assign nG_41_38 = nG_41_40 | (nP_41_40 & nG_39_38);
  assign nP_41_38 = nP_41_40 & nP_39_38;
  assign nG_40_37 = nG_40_39 | (nP_40_39 & nG_38_37);
  assign nP_40_37 = nP_40_39 & nP_38_37;
  assign nG_39_36 = nG_39_38 | (nP_39_38 & nG_37_36);
  assign nP_39_36 = nP_39_38 & nP_37_36;
  assign nG_38_35 = nG_38_37 | (nP_38_37 & nG_36_35);
  assign nP_38_35 = nP_38_37 & nP_36_35;
  assign nG_37_34 = nG_37_36 | (nP_37_36 & nG_35_34);
  assign nP_37_34 = nP_37_36 & nP_35_34;
  assign nG_36_33 = nG_36_35 | (nP_36_35 & nG_34_33);
  assign nP_36_33 = nP_36_35 & nP_34_33;
  assign nG_35_32 = nG_35_34 | (nP_35_34 & nG_33_32);
  assign nP_35_32 = nP_35_34 & nP_33_32;
  assign nG_34_31 = nG_34_33 | (nP_34_33 & nG_32_31);
  assign nP_34_31 = nP_34_33 & nP_32_31;
  assign nG_33_30 = nG_33_32 | (nP_33_32 & nG_31_30);
  assign nP_33_30 = nP_33_32 & nP_31_30;
  assign nG_32_29 = nG_32_31 | (nP_32_31 & nG_30_29);
  assign nP_32_29 = nP_32_31 & nP_30_29;
  assign nG_31_28 = nG_31_30 | (nP_31_30 & nG_29_28);
  assign nP_31_28 = nP_31_30 & nP_29_28;
  assign nG_30_27 = nG_30_29 | (nP_30_29 & nG_28_27);
  assign nP_30_27 = nP_30_29 & nP_28_27;
  assign nG_29_26 = nG_29_28 | (nP_29_28 & nG_27_26);
  assign nP_29_26 = nP_29_28 & nP_27_26;
  assign nG_28_25 = nG_28_27 | (nP_28_27 & nG_26_25);
  assign nP_28_25 = nP_28_27 & nP_26_25;
  assign nG_27_24 = nG_27_26 | (nP_27_26 & nG_25_24);
  assign nP_27_24 = nP_27_26 & nP_25_24;
  assign nG_26_23 = nG_26_25 | (nP_26_25 & nG_24_23);
  assign nP_26_23 = nP_26_25 & nP_24_23;
  assign nG_25_22 = nG_25_24 | (nP_25_24 & nG_23_22);
  assign nP_25_22 = nP_25_24 & nP_23_22;
  assign nG_24_21 = nG_24_23 | (nP_24_23 & nG_22_21);
  assign nP_24_21 = nP_24_23 & nP_22_21;
  assign nG_23_20 = nG_23_22 | (nP_23_22 & nG_21_20);
  assign nP_23_20 = nP_23_22 & nP_21_20;
  assign nG_22_19 = nG_22_21 | (nP_22_21 & nG_20_19);
  assign nP_22_19 = nP_22_21 & nP_20_19;
  assign nG_21_18 = nG_21_20 | (nP_21_20 & nG_19_18);
  assign nP_21_18 = nP_21_20 & nP_19_18;
  assign nG_20_17 = nG_20_19 | (nP_20_19 & nG_18_17);
  assign nP_20_17 = nP_20_19 & nP_18_17;
  assign nG_19_16 = nG_19_18 | (nP_19_18 & nG_17_16);
  assign nP_19_16 = nP_19_18 & nP_17_16;
  assign nG_18_15 = nG_18_17 | (nP_18_17 & nG_16_15);
  assign nP_18_15 = nP_18_17 & nP_16_15;
  assign nG_17_14 = nG_17_16 | (nP_17_16 & nG_15_14);
  assign nP_17_14 = nP_17_16 & nP_15_14;
  assign nG_16_13 = nG_16_15 | (nP_16_15 & nG_14_13);
  assign nP_16_13 = nP_16_15 & nP_14_13;
  assign nG_15_12 = nG_15_14 | (nP_15_14 & nG_13_12);
  assign nP_15_12 = nP_15_14 & nP_13_12;
  assign nG_14_11 = nG_14_13 | (nP_14_13 & nG_12_11);
  assign nP_14_11 = nP_14_13 & nP_12_11;
  assign nG_13_10 = nG_13_12 | (nP_13_12 & nG_11_10);
  assign nP_13_10 = nP_13_12 & nP_11_10;
  assign nG_12_9 = nG_12_11 | (nP_12_11 & nG_10_9);
  assign nP_12_9 = nP_12_11 & nP_10_9;
  assign nG_11_8 = nG_11_10 | (nP_11_10 & nG_9_8);
  assign nP_11_8 = nP_11_10 & nP_9_8;
  assign nG_10_7 = nG_10_9 | (nP_10_9 & nG_8_7);
  assign nP_10_7 = nP_10_9 & nP_8_7;
  assign nG_9_6 = nG_9_8 | (nP_9_8 & nG_7_6);
  assign nP_9_6 = nP_9_8 & nP_7_6;
  assign nG_8_5 = nG_8_7 | (nP_8_7 & nG_6_5);
  assign nP_8_5 = nP_8_7 & nP_6_5;
  assign nG_7_4 = nG_7_6 | (nP_7_6 & nG_5_4);
  assign nP_7_4 = nP_7_6 & nP_5_4;
  assign nG_6_3 = nG_6_5 | (nP_6_5 & nG_4_3);
  assign nP_6_3 = nP_6_5 & nP_4_3;
  assign nG_5_2 = nG_5_4 | (nP_5_4 & nG_3_2);
  assign nP_5_2 = nP_5_4 & nP_3_2;
  assign nG_4_1 = nG_4_3 | (nP_4_3 & nG_2_1);
  assign nP_4_1 = nP_4_3 & nP_2_1;
  assign nG_3_0 = nG_3_2 | (nP_3_2 & nG_1_0);
  assign nP_3_0 = nP_3_2 & nP_1_0;
  assign nG_2_0 = nG_2_1 | (nP_2_1 & nG_0_0);
  assign nP_2_0 = nP_2_1 & nP_0_0;

  assign nG_255_248 = nG_255_252 | (nP_255_252 & nG_251_248);
  assign nP_255_248 = nP_255_252 & nP_251_248;
  assign nG_254_247 = nG_254_251 | (nP_254_251 & nG_250_247);
  assign nP_254_247 = nP_254_251 & nP_250_247;
  assign nG_253_246 = nG_253_250 | (nP_253_250 & nG_249_246);
  assign nP_253_246 = nP_253_250 & nP_249_246;
  assign nG_252_245 = nG_252_249 | (nP_252_249 & nG_248_245);
  assign nP_252_245 = nP_252_249 & nP_248_245;
  assign nG_251_244 = nG_251_248 | (nP_251_248 & nG_247_244);
  assign nP_251_244 = nP_251_248 & nP_247_244;
  assign nG_250_243 = nG_250_247 | (nP_250_247 & nG_246_243);
  assign nP_250_243 = nP_250_247 & nP_246_243;
  assign nG_249_242 = nG_249_246 | (nP_249_246 & nG_245_242);
  assign nP_249_242 = nP_249_246 & nP_245_242;
  assign nG_248_241 = nG_248_245 | (nP_248_245 & nG_244_241);
  assign nP_248_241 = nP_248_245 & nP_244_241;
  assign nG_247_240 = nG_247_244 | (nP_247_244 & nG_243_240);
  assign nP_247_240 = nP_247_244 & nP_243_240;
  assign nG_246_239 = nG_246_243 | (nP_246_243 & nG_242_239);
  assign nP_246_239 = nP_246_243 & nP_242_239;
  assign nG_245_238 = nG_245_242 | (nP_245_242 & nG_241_238);
  assign nP_245_238 = nP_245_242 & nP_241_238;
  assign nG_244_237 = nG_244_241 | (nP_244_241 & nG_240_237);
  assign nP_244_237 = nP_244_241 & nP_240_237;
  assign nG_243_236 = nG_243_240 | (nP_243_240 & nG_239_236);
  assign nP_243_236 = nP_243_240 & nP_239_236;
  assign nG_242_235 = nG_242_239 | (nP_242_239 & nG_238_235);
  assign nP_242_235 = nP_242_239 & nP_238_235;
  assign nG_241_234 = nG_241_238 | (nP_241_238 & nG_237_234);
  assign nP_241_234 = nP_241_238 & nP_237_234;
  assign nG_240_233 = nG_240_237 | (nP_240_237 & nG_236_233);
  assign nP_240_233 = nP_240_237 & nP_236_233;
  assign nG_239_232 = nG_239_236 | (nP_239_236 & nG_235_232);
  assign nP_239_232 = nP_239_236 & nP_235_232;
  assign nG_238_231 = nG_238_235 | (nP_238_235 & nG_234_231);
  assign nP_238_231 = nP_238_235 & nP_234_231;
  assign nG_237_230 = nG_237_234 | (nP_237_234 & nG_233_230);
  assign nP_237_230 = nP_237_234 & nP_233_230;
  assign nG_236_229 = nG_236_233 | (nP_236_233 & nG_232_229);
  assign nP_236_229 = nP_236_233 & nP_232_229;
  assign nG_235_228 = nG_235_232 | (nP_235_232 & nG_231_228);
  assign nP_235_228 = nP_235_232 & nP_231_228;
  assign nG_234_227 = nG_234_231 | (nP_234_231 & nG_230_227);
  assign nP_234_227 = nP_234_231 & nP_230_227;
  assign nG_233_226 = nG_233_230 | (nP_233_230 & nG_229_226);
  assign nP_233_226 = nP_233_230 & nP_229_226;
  assign nG_232_225 = nG_232_229 | (nP_232_229 & nG_228_225);
  assign nP_232_225 = nP_232_229 & nP_228_225;
  assign nG_231_224 = nG_231_228 | (nP_231_228 & nG_227_224);
  assign nP_231_224 = nP_231_228 & nP_227_224;
  assign nG_230_223 = nG_230_227 | (nP_230_227 & nG_226_223);
  assign nP_230_223 = nP_230_227 & nP_226_223;
  assign nG_229_222 = nG_229_226 | (nP_229_226 & nG_225_222);
  assign nP_229_222 = nP_229_226 & nP_225_222;
  assign nG_228_221 = nG_228_225 | (nP_228_225 & nG_224_221);
  assign nP_228_221 = nP_228_225 & nP_224_221;
  assign nG_227_220 = nG_227_224 | (nP_227_224 & nG_223_220);
  assign nP_227_220 = nP_227_224 & nP_223_220;
  assign nG_226_219 = nG_226_223 | (nP_226_223 & nG_222_219);
  assign nP_226_219 = nP_226_223 & nP_222_219;
  assign nG_225_218 = nG_225_222 | (nP_225_222 & nG_221_218);
  assign nP_225_218 = nP_225_222 & nP_221_218;
  assign nG_224_217 = nG_224_221 | (nP_224_221 & nG_220_217);
  assign nP_224_217 = nP_224_221 & nP_220_217;
  assign nG_223_216 = nG_223_220 | (nP_223_220 & nG_219_216);
  assign nP_223_216 = nP_223_220 & nP_219_216;
  assign nG_222_215 = nG_222_219 | (nP_222_219 & nG_218_215);
  assign nP_222_215 = nP_222_219 & nP_218_215;
  assign nG_221_214 = nG_221_218 | (nP_221_218 & nG_217_214);
  assign nP_221_214 = nP_221_218 & nP_217_214;
  assign nG_220_213 = nG_220_217 | (nP_220_217 & nG_216_213);
  assign nP_220_213 = nP_220_217 & nP_216_213;
  assign nG_219_212 = nG_219_216 | (nP_219_216 & nG_215_212);
  assign nP_219_212 = nP_219_216 & nP_215_212;
  assign nG_218_211 = nG_218_215 | (nP_218_215 & nG_214_211);
  assign nP_218_211 = nP_218_215 & nP_214_211;
  assign nG_217_210 = nG_217_214 | (nP_217_214 & nG_213_210);
  assign nP_217_210 = nP_217_214 & nP_213_210;
  assign nG_216_209 = nG_216_213 | (nP_216_213 & nG_212_209);
  assign nP_216_209 = nP_216_213 & nP_212_209;
  assign nG_215_208 = nG_215_212 | (nP_215_212 & nG_211_208);
  assign nP_215_208 = nP_215_212 & nP_211_208;
  assign nG_214_207 = nG_214_211 | (nP_214_211 & nG_210_207);
  assign nP_214_207 = nP_214_211 & nP_210_207;
  assign nG_213_206 = nG_213_210 | (nP_213_210 & nG_209_206);
  assign nP_213_206 = nP_213_210 & nP_209_206;
  assign nG_212_205 = nG_212_209 | (nP_212_209 & nG_208_205);
  assign nP_212_205 = nP_212_209 & nP_208_205;
  assign nG_211_204 = nG_211_208 | (nP_211_208 & nG_207_204);
  assign nP_211_204 = nP_211_208 & nP_207_204;
  assign nG_210_203 = nG_210_207 | (nP_210_207 & nG_206_203);
  assign nP_210_203 = nP_210_207 & nP_206_203;
  assign nG_209_202 = nG_209_206 | (nP_209_206 & nG_205_202);
  assign nP_209_202 = nP_209_206 & nP_205_202;
  assign nG_208_201 = nG_208_205 | (nP_208_205 & nG_204_201);
  assign nP_208_201 = nP_208_205 & nP_204_201;
  assign nG_207_200 = nG_207_204 | (nP_207_204 & nG_203_200);
  assign nP_207_200 = nP_207_204 & nP_203_200;
  assign nG_206_199 = nG_206_203 | (nP_206_203 & nG_202_199);
  assign nP_206_199 = nP_206_203 & nP_202_199;
  assign nG_205_198 = nG_205_202 | (nP_205_202 & nG_201_198);
  assign nP_205_198 = nP_205_202 & nP_201_198;
  assign nG_204_197 = nG_204_201 | (nP_204_201 & nG_200_197);
  assign nP_204_197 = nP_204_201 & nP_200_197;
  assign nG_203_196 = nG_203_200 | (nP_203_200 & nG_199_196);
  assign nP_203_196 = nP_203_200 & nP_199_196;
  assign nG_202_195 = nG_202_199 | (nP_202_199 & nG_198_195);
  assign nP_202_195 = nP_202_199 & nP_198_195;
  assign nG_201_194 = nG_201_198 | (nP_201_198 & nG_197_194);
  assign nP_201_194 = nP_201_198 & nP_197_194;
  assign nG_200_193 = nG_200_197 | (nP_200_197 & nG_196_193);
  assign nP_200_193 = nP_200_197 & nP_196_193;
  assign nG_199_192 = nG_199_196 | (nP_199_196 & nG_195_192);
  assign nP_199_192 = nP_199_196 & nP_195_192;
  assign nG_198_191 = nG_198_195 | (nP_198_195 & nG_194_191);
  assign nP_198_191 = nP_198_195 & nP_194_191;
  assign nG_197_190 = nG_197_194 | (nP_197_194 & nG_193_190);
  assign nP_197_190 = nP_197_194 & nP_193_190;
  assign nG_196_189 = nG_196_193 | (nP_196_193 & nG_192_189);
  assign nP_196_189 = nP_196_193 & nP_192_189;
  assign nG_195_188 = nG_195_192 | (nP_195_192 & nG_191_188);
  assign nP_195_188 = nP_195_192 & nP_191_188;
  assign nG_194_187 = nG_194_191 | (nP_194_191 & nG_190_187);
  assign nP_194_187 = nP_194_191 & nP_190_187;
  assign nG_193_186 = nG_193_190 | (nP_193_190 & nG_189_186);
  assign nP_193_186 = nP_193_190 & nP_189_186;
  assign nG_192_185 = nG_192_189 | (nP_192_189 & nG_188_185);
  assign nP_192_185 = nP_192_189 & nP_188_185;
  assign nG_191_184 = nG_191_188 | (nP_191_188 & nG_187_184);
  assign nP_191_184 = nP_191_188 & nP_187_184;
  assign nG_190_183 = nG_190_187 | (nP_190_187 & nG_186_183);
  assign nP_190_183 = nP_190_187 & nP_186_183;
  assign nG_189_182 = nG_189_186 | (nP_189_186 & nG_185_182);
  assign nP_189_182 = nP_189_186 & nP_185_182;
  assign nG_188_181 = nG_188_185 | (nP_188_185 & nG_184_181);
  assign nP_188_181 = nP_188_185 & nP_184_181;
  assign nG_187_180 = nG_187_184 | (nP_187_184 & nG_183_180);
  assign nP_187_180 = nP_187_184 & nP_183_180;
  assign nG_186_179 = nG_186_183 | (nP_186_183 & nG_182_179);
  assign nP_186_179 = nP_186_183 & nP_182_179;
  assign nG_185_178 = nG_185_182 | (nP_185_182 & nG_181_178);
  assign nP_185_178 = nP_185_182 & nP_181_178;
  assign nG_184_177 = nG_184_181 | (nP_184_181 & nG_180_177);
  assign nP_184_177 = nP_184_181 & nP_180_177;
  assign nG_183_176 = nG_183_180 | (nP_183_180 & nG_179_176);
  assign nP_183_176 = nP_183_180 & nP_179_176;
  assign nG_182_175 = nG_182_179 | (nP_182_179 & nG_178_175);
  assign nP_182_175 = nP_182_179 & nP_178_175;
  assign nG_181_174 = nG_181_178 | (nP_181_178 & nG_177_174);
  assign nP_181_174 = nP_181_178 & nP_177_174;
  assign nG_180_173 = nG_180_177 | (nP_180_177 & nG_176_173);
  assign nP_180_173 = nP_180_177 & nP_176_173;
  assign nG_179_172 = nG_179_176 | (nP_179_176 & nG_175_172);
  assign nP_179_172 = nP_179_176 & nP_175_172;
  assign nG_178_171 = nG_178_175 | (nP_178_175 & nG_174_171);
  assign nP_178_171 = nP_178_175 & nP_174_171;
  assign nG_177_170 = nG_177_174 | (nP_177_174 & nG_173_170);
  assign nP_177_170 = nP_177_174 & nP_173_170;
  assign nG_176_169 = nG_176_173 | (nP_176_173 & nG_172_169);
  assign nP_176_169 = nP_176_173 & nP_172_169;
  assign nG_175_168 = nG_175_172 | (nP_175_172 & nG_171_168);
  assign nP_175_168 = nP_175_172 & nP_171_168;
  assign nG_174_167 = nG_174_171 | (nP_174_171 & nG_170_167);
  assign nP_174_167 = nP_174_171 & nP_170_167;
  assign nG_173_166 = nG_173_170 | (nP_173_170 & nG_169_166);
  assign nP_173_166 = nP_173_170 & nP_169_166;
  assign nG_172_165 = nG_172_169 | (nP_172_169 & nG_168_165);
  assign nP_172_165 = nP_172_169 & nP_168_165;
  assign nG_171_164 = nG_171_168 | (nP_171_168 & nG_167_164);
  assign nP_171_164 = nP_171_168 & nP_167_164;
  assign nG_170_163 = nG_170_167 | (nP_170_167 & nG_166_163);
  assign nP_170_163 = nP_170_167 & nP_166_163;
  assign nG_169_162 = nG_169_166 | (nP_169_166 & nG_165_162);
  assign nP_169_162 = nP_169_166 & nP_165_162;
  assign nG_168_161 = nG_168_165 | (nP_168_165 & nG_164_161);
  assign nP_168_161 = nP_168_165 & nP_164_161;
  assign nG_167_160 = nG_167_164 | (nP_167_164 & nG_163_160);
  assign nP_167_160 = nP_167_164 & nP_163_160;
  assign nG_166_159 = nG_166_163 | (nP_166_163 & nG_162_159);
  assign nP_166_159 = nP_166_163 & nP_162_159;
  assign nG_165_158 = nG_165_162 | (nP_165_162 & nG_161_158);
  assign nP_165_158 = nP_165_162 & nP_161_158;
  assign nG_164_157 = nG_164_161 | (nP_164_161 & nG_160_157);
  assign nP_164_157 = nP_164_161 & nP_160_157;
  assign nG_163_156 = nG_163_160 | (nP_163_160 & nG_159_156);
  assign nP_163_156 = nP_163_160 & nP_159_156;
  assign nG_162_155 = nG_162_159 | (nP_162_159 & nG_158_155);
  assign nP_162_155 = nP_162_159 & nP_158_155;
  assign nG_161_154 = nG_161_158 | (nP_161_158 & nG_157_154);
  assign nP_161_154 = nP_161_158 & nP_157_154;
  assign nG_160_153 = nG_160_157 | (nP_160_157 & nG_156_153);
  assign nP_160_153 = nP_160_157 & nP_156_153;
  assign nG_159_152 = nG_159_156 | (nP_159_156 & nG_155_152);
  assign nP_159_152 = nP_159_156 & nP_155_152;
  assign nG_158_151 = nG_158_155 | (nP_158_155 & nG_154_151);
  assign nP_158_151 = nP_158_155 & nP_154_151;
  assign nG_157_150 = nG_157_154 | (nP_157_154 & nG_153_150);
  assign nP_157_150 = nP_157_154 & nP_153_150;
  assign nG_156_149 = nG_156_153 | (nP_156_153 & nG_152_149);
  assign nP_156_149 = nP_156_153 & nP_152_149;
  assign nG_155_148 = nG_155_152 | (nP_155_152 & nG_151_148);
  assign nP_155_148 = nP_155_152 & nP_151_148;
  assign nG_154_147 = nG_154_151 | (nP_154_151 & nG_150_147);
  assign nP_154_147 = nP_154_151 & nP_150_147;
  assign nG_153_146 = nG_153_150 | (nP_153_150 & nG_149_146);
  assign nP_153_146 = nP_153_150 & nP_149_146;
  assign nG_152_145 = nG_152_149 | (nP_152_149 & nG_148_145);
  assign nP_152_145 = nP_152_149 & nP_148_145;
  assign nG_151_144 = nG_151_148 | (nP_151_148 & nG_147_144);
  assign nP_151_144 = nP_151_148 & nP_147_144;
  assign nG_150_143 = nG_150_147 | (nP_150_147 & nG_146_143);
  assign nP_150_143 = nP_150_147 & nP_146_143;
  assign nG_149_142 = nG_149_146 | (nP_149_146 & nG_145_142);
  assign nP_149_142 = nP_149_146 & nP_145_142;
  assign nG_148_141 = nG_148_145 | (nP_148_145 & nG_144_141);
  assign nP_148_141 = nP_148_145 & nP_144_141;
  assign nG_147_140 = nG_147_144 | (nP_147_144 & nG_143_140);
  assign nP_147_140 = nP_147_144 & nP_143_140;
  assign nG_146_139 = nG_146_143 | (nP_146_143 & nG_142_139);
  assign nP_146_139 = nP_146_143 & nP_142_139;
  assign nG_145_138 = nG_145_142 | (nP_145_142 & nG_141_138);
  assign nP_145_138 = nP_145_142 & nP_141_138;
  assign nG_144_137 = nG_144_141 | (nP_144_141 & nG_140_137);
  assign nP_144_137 = nP_144_141 & nP_140_137;
  assign nG_143_136 = nG_143_140 | (nP_143_140 & nG_139_136);
  assign nP_143_136 = nP_143_140 & nP_139_136;
  assign nG_142_135 = nG_142_139 | (nP_142_139 & nG_138_135);
  assign nP_142_135 = nP_142_139 & nP_138_135;
  assign nG_141_134 = nG_141_138 | (nP_141_138 & nG_137_134);
  assign nP_141_134 = nP_141_138 & nP_137_134;
  assign nG_140_133 = nG_140_137 | (nP_140_137 & nG_136_133);
  assign nP_140_133 = nP_140_137 & nP_136_133;
  assign nG_139_132 = nG_139_136 | (nP_139_136 & nG_135_132);
  assign nP_139_132 = nP_139_136 & nP_135_132;
  assign nG_138_131 = nG_138_135 | (nP_138_135 & nG_134_131);
  assign nP_138_131 = nP_138_135 & nP_134_131;
  assign nG_137_130 = nG_137_134 | (nP_137_134 & nG_133_130);
  assign nP_137_130 = nP_137_134 & nP_133_130;
  assign nG_136_129 = nG_136_133 | (nP_136_133 & nG_132_129);
  assign nP_136_129 = nP_136_133 & nP_132_129;
  assign nG_135_128 = nG_135_132 | (nP_135_132 & nG_131_128);
  assign nP_135_128 = nP_135_132 & nP_131_128;
  assign nG_134_127 = nG_134_131 | (nP_134_131 & nG_130_127);
  assign nP_134_127 = nP_134_131 & nP_130_127;
  assign nG_133_126 = nG_133_130 | (nP_133_130 & nG_129_126);
  assign nP_133_126 = nP_133_130 & nP_129_126;
  assign nG_132_125 = nG_132_129 | (nP_132_129 & nG_128_125);
  assign nP_132_125 = nP_132_129 & nP_128_125;
  assign nG_131_124 = nG_131_128 | (nP_131_128 & nG_127_124);
  assign nP_131_124 = nP_131_128 & nP_127_124;
  assign nG_130_123 = nG_130_127 | (nP_130_127 & nG_126_123);
  assign nP_130_123 = nP_130_127 & nP_126_123;
  assign nG_129_122 = nG_129_126 | (nP_129_126 & nG_125_122);
  assign nP_129_122 = nP_129_126 & nP_125_122;
  assign nG_128_121 = nG_128_125 | (nP_128_125 & nG_124_121);
  assign nP_128_121 = nP_128_125 & nP_124_121;
  assign nG_127_120 = nG_127_124 | (nP_127_124 & nG_123_120);
  assign nP_127_120 = nP_127_124 & nP_123_120;
  assign nG_126_119 = nG_126_123 | (nP_126_123 & nG_122_119);
  assign nP_126_119 = nP_126_123 & nP_122_119;
  assign nG_125_118 = nG_125_122 | (nP_125_122 & nG_121_118);
  assign nP_125_118 = nP_125_122 & nP_121_118;
  assign nG_124_117 = nG_124_121 | (nP_124_121 & nG_120_117);
  assign nP_124_117 = nP_124_121 & nP_120_117;
  assign nG_123_116 = nG_123_120 | (nP_123_120 & nG_119_116);
  assign nP_123_116 = nP_123_120 & nP_119_116;
  assign nG_122_115 = nG_122_119 | (nP_122_119 & nG_118_115);
  assign nP_122_115 = nP_122_119 & nP_118_115;
  assign nG_121_114 = nG_121_118 | (nP_121_118 & nG_117_114);
  assign nP_121_114 = nP_121_118 & nP_117_114;
  assign nG_120_113 = nG_120_117 | (nP_120_117 & nG_116_113);
  assign nP_120_113 = nP_120_117 & nP_116_113;
  assign nG_119_112 = nG_119_116 | (nP_119_116 & nG_115_112);
  assign nP_119_112 = nP_119_116 & nP_115_112;
  assign nG_118_111 = nG_118_115 | (nP_118_115 & nG_114_111);
  assign nP_118_111 = nP_118_115 & nP_114_111;
  assign nG_117_110 = nG_117_114 | (nP_117_114 & nG_113_110);
  assign nP_117_110 = nP_117_114 & nP_113_110;
  assign nG_116_109 = nG_116_113 | (nP_116_113 & nG_112_109);
  assign nP_116_109 = nP_116_113 & nP_112_109;
  assign nG_115_108 = nG_115_112 | (nP_115_112 & nG_111_108);
  assign nP_115_108 = nP_115_112 & nP_111_108;
  assign nG_114_107 = nG_114_111 | (nP_114_111 & nG_110_107);
  assign nP_114_107 = nP_114_111 & nP_110_107;
  assign nG_113_106 = nG_113_110 | (nP_113_110 & nG_109_106);
  assign nP_113_106 = nP_113_110 & nP_109_106;
  assign nG_112_105 = nG_112_109 | (nP_112_109 & nG_108_105);
  assign nP_112_105 = nP_112_109 & nP_108_105;
  assign nG_111_104 = nG_111_108 | (nP_111_108 & nG_107_104);
  assign nP_111_104 = nP_111_108 & nP_107_104;
  assign nG_110_103 = nG_110_107 | (nP_110_107 & nG_106_103);
  assign nP_110_103 = nP_110_107 & nP_106_103;
  assign nG_109_102 = nG_109_106 | (nP_109_106 & nG_105_102);
  assign nP_109_102 = nP_109_106 & nP_105_102;
  assign nG_108_101 = nG_108_105 | (nP_108_105 & nG_104_101);
  assign nP_108_101 = nP_108_105 & nP_104_101;
  assign nG_107_100 = nG_107_104 | (nP_107_104 & nG_103_100);
  assign nP_107_100 = nP_107_104 & nP_103_100;
  assign nG_106_99 = nG_106_103 | (nP_106_103 & nG_102_99);
  assign nP_106_99 = nP_106_103 & nP_102_99;
  assign nG_105_98 = nG_105_102 | (nP_105_102 & nG_101_98);
  assign nP_105_98 = nP_105_102 & nP_101_98;
  assign nG_104_97 = nG_104_101 | (nP_104_101 & nG_100_97);
  assign nP_104_97 = nP_104_101 & nP_100_97;
  assign nG_103_96 = nG_103_100 | (nP_103_100 & nG_99_96);
  assign nP_103_96 = nP_103_100 & nP_99_96;
  assign nG_102_95 = nG_102_99 | (nP_102_99 & nG_98_95);
  assign nP_102_95 = nP_102_99 & nP_98_95;
  assign nG_101_94 = nG_101_98 | (nP_101_98 & nG_97_94);
  assign nP_101_94 = nP_101_98 & nP_97_94;
  assign nG_100_93 = nG_100_97 | (nP_100_97 & nG_96_93);
  assign nP_100_93 = nP_100_97 & nP_96_93;
  assign nG_99_92 = nG_99_96 | (nP_99_96 & nG_95_92);
  assign nP_99_92 = nP_99_96 & nP_95_92;
  assign nG_98_91 = nG_98_95 | (nP_98_95 & nG_94_91);
  assign nP_98_91 = nP_98_95 & nP_94_91;
  assign nG_97_90 = nG_97_94 | (nP_97_94 & nG_93_90);
  assign nP_97_90 = nP_97_94 & nP_93_90;
  assign nG_96_89 = nG_96_93 | (nP_96_93 & nG_92_89);
  assign nP_96_89 = nP_96_93 & nP_92_89;
  assign nG_95_88 = nG_95_92 | (nP_95_92 & nG_91_88);
  assign nP_95_88 = nP_95_92 & nP_91_88;
  assign nG_94_87 = nG_94_91 | (nP_94_91 & nG_90_87);
  assign nP_94_87 = nP_94_91 & nP_90_87;
  assign nG_93_86 = nG_93_90 | (nP_93_90 & nG_89_86);
  assign nP_93_86 = nP_93_90 & nP_89_86;
  assign nG_92_85 = nG_92_89 | (nP_92_89 & nG_88_85);
  assign nP_92_85 = nP_92_89 & nP_88_85;
  assign nG_91_84 = nG_91_88 | (nP_91_88 & nG_87_84);
  assign nP_91_84 = nP_91_88 & nP_87_84;
  assign nG_90_83 = nG_90_87 | (nP_90_87 & nG_86_83);
  assign nP_90_83 = nP_90_87 & nP_86_83;
  assign nG_89_82 = nG_89_86 | (nP_89_86 & nG_85_82);
  assign nP_89_82 = nP_89_86 & nP_85_82;
  assign nG_88_81 = nG_88_85 | (nP_88_85 & nG_84_81);
  assign nP_88_81 = nP_88_85 & nP_84_81;
  assign nG_87_80 = nG_87_84 | (nP_87_84 & nG_83_80);
  assign nP_87_80 = nP_87_84 & nP_83_80;
  assign nG_86_79 = nG_86_83 | (nP_86_83 & nG_82_79);
  assign nP_86_79 = nP_86_83 & nP_82_79;
  assign nG_85_78 = nG_85_82 | (nP_85_82 & nG_81_78);
  assign nP_85_78 = nP_85_82 & nP_81_78;
  assign nG_84_77 = nG_84_81 | (nP_84_81 & nG_80_77);
  assign nP_84_77 = nP_84_81 & nP_80_77;
  assign nG_83_76 = nG_83_80 | (nP_83_80 & nG_79_76);
  assign nP_83_76 = nP_83_80 & nP_79_76;
  assign nG_82_75 = nG_82_79 | (nP_82_79 & nG_78_75);
  assign nP_82_75 = nP_82_79 & nP_78_75;
  assign nG_81_74 = nG_81_78 | (nP_81_78 & nG_77_74);
  assign nP_81_74 = nP_81_78 & nP_77_74;
  assign nG_80_73 = nG_80_77 | (nP_80_77 & nG_76_73);
  assign nP_80_73 = nP_80_77 & nP_76_73;
  assign nG_79_72 = nG_79_76 | (nP_79_76 & nG_75_72);
  assign nP_79_72 = nP_79_76 & nP_75_72;
  assign nG_78_71 = nG_78_75 | (nP_78_75 & nG_74_71);
  assign nP_78_71 = nP_78_75 & nP_74_71;
  assign nG_77_70 = nG_77_74 | (nP_77_74 & nG_73_70);
  assign nP_77_70 = nP_77_74 & nP_73_70;
  assign nG_76_69 = nG_76_73 | (nP_76_73 & nG_72_69);
  assign nP_76_69 = nP_76_73 & nP_72_69;
  assign nG_75_68 = nG_75_72 | (nP_75_72 & nG_71_68);
  assign nP_75_68 = nP_75_72 & nP_71_68;
  assign nG_74_67 = nG_74_71 | (nP_74_71 & nG_70_67);
  assign nP_74_67 = nP_74_71 & nP_70_67;
  assign nG_73_66 = nG_73_70 | (nP_73_70 & nG_69_66);
  assign nP_73_66 = nP_73_70 & nP_69_66;
  assign nG_72_65 = nG_72_69 | (nP_72_69 & nG_68_65);
  assign nP_72_65 = nP_72_69 & nP_68_65;
  assign nG_71_64 = nG_71_68 | (nP_71_68 & nG_67_64);
  assign nP_71_64 = nP_71_68 & nP_67_64;
  assign nG_70_63 = nG_70_67 | (nP_70_67 & nG_66_63);
  assign nP_70_63 = nP_70_67 & nP_66_63;
  assign nG_69_62 = nG_69_66 | (nP_69_66 & nG_65_62);
  assign nP_69_62 = nP_69_66 & nP_65_62;
  assign nG_68_61 = nG_68_65 | (nP_68_65 & nG_64_61);
  assign nP_68_61 = nP_68_65 & nP_64_61;
  assign nG_67_60 = nG_67_64 | (nP_67_64 & nG_63_60);
  assign nP_67_60 = nP_67_64 & nP_63_60;
  assign nG_66_59 = nG_66_63 | (nP_66_63 & nG_62_59);
  assign nP_66_59 = nP_66_63 & nP_62_59;
  assign nG_65_58 = nG_65_62 | (nP_65_62 & nG_61_58);
  assign nP_65_58 = nP_65_62 & nP_61_58;
  assign nG_64_57 = nG_64_61 | (nP_64_61 & nG_60_57);
  assign nP_64_57 = nP_64_61 & nP_60_57;
  assign nG_63_56 = nG_63_60 | (nP_63_60 & nG_59_56);
  assign nP_63_56 = nP_63_60 & nP_59_56;
  assign nG_62_55 = nG_62_59 | (nP_62_59 & nG_58_55);
  assign nP_62_55 = nP_62_59 & nP_58_55;
  assign nG_61_54 = nG_61_58 | (nP_61_58 & nG_57_54);
  assign nP_61_54 = nP_61_58 & nP_57_54;
  assign nG_60_53 = nG_60_57 | (nP_60_57 & nG_56_53);
  assign nP_60_53 = nP_60_57 & nP_56_53;
  assign nG_59_52 = nG_59_56 | (nP_59_56 & nG_55_52);
  assign nP_59_52 = nP_59_56 & nP_55_52;
  assign nG_58_51 = nG_58_55 | (nP_58_55 & nG_54_51);
  assign nP_58_51 = nP_58_55 & nP_54_51;
  assign nG_57_50 = nG_57_54 | (nP_57_54 & nG_53_50);
  assign nP_57_50 = nP_57_54 & nP_53_50;
  assign nG_56_49 = nG_56_53 | (nP_56_53 & nG_52_49);
  assign nP_56_49 = nP_56_53 & nP_52_49;
  assign nG_55_48 = nG_55_52 | (nP_55_52 & nG_51_48);
  assign nP_55_48 = nP_55_52 & nP_51_48;
  assign nG_54_47 = nG_54_51 | (nP_54_51 & nG_50_47);
  assign nP_54_47 = nP_54_51 & nP_50_47;
  assign nG_53_46 = nG_53_50 | (nP_53_50 & nG_49_46);
  assign nP_53_46 = nP_53_50 & nP_49_46;
  assign nG_52_45 = nG_52_49 | (nP_52_49 & nG_48_45);
  assign nP_52_45 = nP_52_49 & nP_48_45;
  assign nG_51_44 = nG_51_48 | (nP_51_48 & nG_47_44);
  assign nP_51_44 = nP_51_48 & nP_47_44;
  assign nG_50_43 = nG_50_47 | (nP_50_47 & nG_46_43);
  assign nP_50_43 = nP_50_47 & nP_46_43;
  assign nG_49_42 = nG_49_46 | (nP_49_46 & nG_45_42);
  assign nP_49_42 = nP_49_46 & nP_45_42;
  assign nG_48_41 = nG_48_45 | (nP_48_45 & nG_44_41);
  assign nP_48_41 = nP_48_45 & nP_44_41;
  assign nG_47_40 = nG_47_44 | (nP_47_44 & nG_43_40);
  assign nP_47_40 = nP_47_44 & nP_43_40;
  assign nG_46_39 = nG_46_43 | (nP_46_43 & nG_42_39);
  assign nP_46_39 = nP_46_43 & nP_42_39;
  assign nG_45_38 = nG_45_42 | (nP_45_42 & nG_41_38);
  assign nP_45_38 = nP_45_42 & nP_41_38;
  assign nG_44_37 = nG_44_41 | (nP_44_41 & nG_40_37);
  assign nP_44_37 = nP_44_41 & nP_40_37;
  assign nG_43_36 = nG_43_40 | (nP_43_40 & nG_39_36);
  assign nP_43_36 = nP_43_40 & nP_39_36;
  assign nG_42_35 = nG_42_39 | (nP_42_39 & nG_38_35);
  assign nP_42_35 = nP_42_39 & nP_38_35;
  assign nG_41_34 = nG_41_38 | (nP_41_38 & nG_37_34);
  assign nP_41_34 = nP_41_38 & nP_37_34;
  assign nG_40_33 = nG_40_37 | (nP_40_37 & nG_36_33);
  assign nP_40_33 = nP_40_37 & nP_36_33;
  assign nG_39_32 = nG_39_36 | (nP_39_36 & nG_35_32);
  assign nP_39_32 = nP_39_36 & nP_35_32;
  assign nG_38_31 = nG_38_35 | (nP_38_35 & nG_34_31);
  assign nP_38_31 = nP_38_35 & nP_34_31;
  assign nG_37_30 = nG_37_34 | (nP_37_34 & nG_33_30);
  assign nP_37_30 = nP_37_34 & nP_33_30;
  assign nG_36_29 = nG_36_33 | (nP_36_33 & nG_32_29);
  assign nP_36_29 = nP_36_33 & nP_32_29;
  assign nG_35_28 = nG_35_32 | (nP_35_32 & nG_31_28);
  assign nP_35_28 = nP_35_32 & nP_31_28;
  assign nG_34_27 = nG_34_31 | (nP_34_31 & nG_30_27);
  assign nP_34_27 = nP_34_31 & nP_30_27;
  assign nG_33_26 = nG_33_30 | (nP_33_30 & nG_29_26);
  assign nP_33_26 = nP_33_30 & nP_29_26;
  assign nG_32_25 = nG_32_29 | (nP_32_29 & nG_28_25);
  assign nP_32_25 = nP_32_29 & nP_28_25;
  assign nG_31_24 = nG_31_28 | (nP_31_28 & nG_27_24);
  assign nP_31_24 = nP_31_28 & nP_27_24;
  assign nG_30_23 = nG_30_27 | (nP_30_27 & nG_26_23);
  assign nP_30_23 = nP_30_27 & nP_26_23;
  assign nG_29_22 = nG_29_26 | (nP_29_26 & nG_25_22);
  assign nP_29_22 = nP_29_26 & nP_25_22;
  assign nG_28_21 = nG_28_25 | (nP_28_25 & nG_24_21);
  assign nP_28_21 = nP_28_25 & nP_24_21;
  assign nG_27_20 = nG_27_24 | (nP_27_24 & nG_23_20);
  assign nP_27_20 = nP_27_24 & nP_23_20;
  assign nG_26_19 = nG_26_23 | (nP_26_23 & nG_22_19);
  assign nP_26_19 = nP_26_23 & nP_22_19;
  assign nG_25_18 = nG_25_22 | (nP_25_22 & nG_21_18);
  assign nP_25_18 = nP_25_22 & nP_21_18;
  assign nG_24_17 = nG_24_21 | (nP_24_21 & nG_20_17);
  assign nP_24_17 = nP_24_21 & nP_20_17;
  assign nG_23_16 = nG_23_20 | (nP_23_20 & nG_19_16);
  assign nP_23_16 = nP_23_20 & nP_19_16;
  assign nG_22_15 = nG_22_19 | (nP_22_19 & nG_18_15);
  assign nP_22_15 = nP_22_19 & nP_18_15;
  assign nG_21_14 = nG_21_18 | (nP_21_18 & nG_17_14);
  assign nP_21_14 = nP_21_18 & nP_17_14;
  assign nG_20_13 = nG_20_17 | (nP_20_17 & nG_16_13);
  assign nP_20_13 = nP_20_17 & nP_16_13;
  assign nG_19_12 = nG_19_16 | (nP_19_16 & nG_15_12);
  assign nP_19_12 = nP_19_16 & nP_15_12;
  assign nG_18_11 = nG_18_15 | (nP_18_15 & nG_14_11);
  assign nP_18_11 = nP_18_15 & nP_14_11;
  assign nG_17_10 = nG_17_14 | (nP_17_14 & nG_13_10);
  assign nP_17_10 = nP_17_14 & nP_13_10;
  assign nG_16_9 = nG_16_13 | (nP_16_13 & nG_12_9);
  assign nP_16_9 = nP_16_13 & nP_12_9;
  assign nG_15_8 = nG_15_12 | (nP_15_12 & nG_11_8);
  assign nP_15_8 = nP_15_12 & nP_11_8;
  assign nG_14_7 = nG_14_11 | (nP_14_11 & nG_10_7);
  assign nP_14_7 = nP_14_11 & nP_10_7;
  assign nG_13_6 = nG_13_10 | (nP_13_10 & nG_9_6);
  assign nP_13_6 = nP_13_10 & nP_9_6;
  assign nG_12_5 = nG_12_9 | (nP_12_9 & nG_8_5);
  assign nP_12_5 = nP_12_9 & nP_8_5;
  assign nG_11_4 = nG_11_8 | (nP_11_8 & nG_7_4);
  assign nP_11_4 = nP_11_8 & nP_7_4;
  assign nG_10_3 = nG_10_7 | (nP_10_7 & nG_6_3);
  assign nP_10_3 = nP_10_7 & nP_6_3;
  assign nG_9_2 = nG_9_6 | (nP_9_6 & nG_5_2);
  assign nP_9_2 = nP_9_6 & nP_5_2;
  assign nG_8_1 = nG_8_5 | (nP_8_5 & nG_4_1);
  assign nP_8_1 = nP_8_5 & nP_4_1;
  assign nG_7_0 = nG_7_4 | (nP_7_4 & nG_3_0);
  assign nP_7_0 = nP_7_4 & nP_3_0;
  assign nG_6_0 = nG_6_3 | (nP_6_3 & nG_2_0);
  assign nP_6_0 = nP_6_3 & nP_2_0;
  assign nG_5_0 = nG_5_2 | (nP_5_2 & nG_1_0);
  assign nP_5_0 = nP_5_2 & nP_1_0;
  assign nG_4_0 = nG_4_1 | (nP_4_1 & nG_0_0);
  assign nP_4_0 = nP_4_1 & nP_0_0;

  assign nG_255_240 = nG_255_248 | (nP_255_248 & nG_247_240);
  assign nP_255_240 = nP_255_248 & nP_247_240;
  assign nG_254_239 = nG_254_247 | (nP_254_247 & nG_246_239);
  assign nP_254_239 = nP_254_247 & nP_246_239;
  assign nG_253_238 = nG_253_246 | (nP_253_246 & nG_245_238);
  assign nP_253_238 = nP_253_246 & nP_245_238;
  assign nG_252_237 = nG_252_245 | (nP_252_245 & nG_244_237);
  assign nP_252_237 = nP_252_245 & nP_244_237;
  assign nG_251_236 = nG_251_244 | (nP_251_244 & nG_243_236);
  assign nP_251_236 = nP_251_244 & nP_243_236;
  assign nG_250_235 = nG_250_243 | (nP_250_243 & nG_242_235);
  assign nP_250_235 = nP_250_243 & nP_242_235;
  assign nG_249_234 = nG_249_242 | (nP_249_242 & nG_241_234);
  assign nP_249_234 = nP_249_242 & nP_241_234;
  assign nG_248_233 = nG_248_241 | (nP_248_241 & nG_240_233);
  assign nP_248_233 = nP_248_241 & nP_240_233;
  assign nG_247_232 = nG_247_240 | (nP_247_240 & nG_239_232);
  assign nP_247_232 = nP_247_240 & nP_239_232;
  assign nG_246_231 = nG_246_239 | (nP_246_239 & nG_238_231);
  assign nP_246_231 = nP_246_239 & nP_238_231;
  assign nG_245_230 = nG_245_238 | (nP_245_238 & nG_237_230);
  assign nP_245_230 = nP_245_238 & nP_237_230;
  assign nG_244_229 = nG_244_237 | (nP_244_237 & nG_236_229);
  assign nP_244_229 = nP_244_237 & nP_236_229;
  assign nG_243_228 = nG_243_236 | (nP_243_236 & nG_235_228);
  assign nP_243_228 = nP_243_236 & nP_235_228;
  assign nG_242_227 = nG_242_235 | (nP_242_235 & nG_234_227);
  assign nP_242_227 = nP_242_235 & nP_234_227;
  assign nG_241_226 = nG_241_234 | (nP_241_234 & nG_233_226);
  assign nP_241_226 = nP_241_234 & nP_233_226;
  assign nG_240_225 = nG_240_233 | (nP_240_233 & nG_232_225);
  assign nP_240_225 = nP_240_233 & nP_232_225;
  assign nG_239_224 = nG_239_232 | (nP_239_232 & nG_231_224);
  assign nP_239_224 = nP_239_232 & nP_231_224;
  assign nG_238_223 = nG_238_231 | (nP_238_231 & nG_230_223);
  assign nP_238_223 = nP_238_231 & nP_230_223;
  assign nG_237_222 = nG_237_230 | (nP_237_230 & nG_229_222);
  assign nP_237_222 = nP_237_230 & nP_229_222;
  assign nG_236_221 = nG_236_229 | (nP_236_229 & nG_228_221);
  assign nP_236_221 = nP_236_229 & nP_228_221;
  assign nG_235_220 = nG_235_228 | (nP_235_228 & nG_227_220);
  assign nP_235_220 = nP_235_228 & nP_227_220;
  assign nG_234_219 = nG_234_227 | (nP_234_227 & nG_226_219);
  assign nP_234_219 = nP_234_227 & nP_226_219;
  assign nG_233_218 = nG_233_226 | (nP_233_226 & nG_225_218);
  assign nP_233_218 = nP_233_226 & nP_225_218;
  assign nG_232_217 = nG_232_225 | (nP_232_225 & nG_224_217);
  assign nP_232_217 = nP_232_225 & nP_224_217;
  assign nG_231_216 = nG_231_224 | (nP_231_224 & nG_223_216);
  assign nP_231_216 = nP_231_224 & nP_223_216;
  assign nG_230_215 = nG_230_223 | (nP_230_223 & nG_222_215);
  assign nP_230_215 = nP_230_223 & nP_222_215;
  assign nG_229_214 = nG_229_222 | (nP_229_222 & nG_221_214);
  assign nP_229_214 = nP_229_222 & nP_221_214;
  assign nG_228_213 = nG_228_221 | (nP_228_221 & nG_220_213);
  assign nP_228_213 = nP_228_221 & nP_220_213;
  assign nG_227_212 = nG_227_220 | (nP_227_220 & nG_219_212);
  assign nP_227_212 = nP_227_220 & nP_219_212;
  assign nG_226_211 = nG_226_219 | (nP_226_219 & nG_218_211);
  assign nP_226_211 = nP_226_219 & nP_218_211;
  assign nG_225_210 = nG_225_218 | (nP_225_218 & nG_217_210);
  assign nP_225_210 = nP_225_218 & nP_217_210;
  assign nG_224_209 = nG_224_217 | (nP_224_217 & nG_216_209);
  assign nP_224_209 = nP_224_217 & nP_216_209;
  assign nG_223_208 = nG_223_216 | (nP_223_216 & nG_215_208);
  assign nP_223_208 = nP_223_216 & nP_215_208;
  assign nG_222_207 = nG_222_215 | (nP_222_215 & nG_214_207);
  assign nP_222_207 = nP_222_215 & nP_214_207;
  assign nG_221_206 = nG_221_214 | (nP_221_214 & nG_213_206);
  assign nP_221_206 = nP_221_214 & nP_213_206;
  assign nG_220_205 = nG_220_213 | (nP_220_213 & nG_212_205);
  assign nP_220_205 = nP_220_213 & nP_212_205;
  assign nG_219_204 = nG_219_212 | (nP_219_212 & nG_211_204);
  assign nP_219_204 = nP_219_212 & nP_211_204;
  assign nG_218_203 = nG_218_211 | (nP_218_211 & nG_210_203);
  assign nP_218_203 = nP_218_211 & nP_210_203;
  assign nG_217_202 = nG_217_210 | (nP_217_210 & nG_209_202);
  assign nP_217_202 = nP_217_210 & nP_209_202;
  assign nG_216_201 = nG_216_209 | (nP_216_209 & nG_208_201);
  assign nP_216_201 = nP_216_209 & nP_208_201;
  assign nG_215_200 = nG_215_208 | (nP_215_208 & nG_207_200);
  assign nP_215_200 = nP_215_208 & nP_207_200;
  assign nG_214_199 = nG_214_207 | (nP_214_207 & nG_206_199);
  assign nP_214_199 = nP_214_207 & nP_206_199;
  assign nG_213_198 = nG_213_206 | (nP_213_206 & nG_205_198);
  assign nP_213_198 = nP_213_206 & nP_205_198;
  assign nG_212_197 = nG_212_205 | (nP_212_205 & nG_204_197);
  assign nP_212_197 = nP_212_205 & nP_204_197;
  assign nG_211_196 = nG_211_204 | (nP_211_204 & nG_203_196);
  assign nP_211_196 = nP_211_204 & nP_203_196;
  assign nG_210_195 = nG_210_203 | (nP_210_203 & nG_202_195);
  assign nP_210_195 = nP_210_203 & nP_202_195;
  assign nG_209_194 = nG_209_202 | (nP_209_202 & nG_201_194);
  assign nP_209_194 = nP_209_202 & nP_201_194;
  assign nG_208_193 = nG_208_201 | (nP_208_201 & nG_200_193);
  assign nP_208_193 = nP_208_201 & nP_200_193;
  assign nG_207_192 = nG_207_200 | (nP_207_200 & nG_199_192);
  assign nP_207_192 = nP_207_200 & nP_199_192;
  assign nG_206_191 = nG_206_199 | (nP_206_199 & nG_198_191);
  assign nP_206_191 = nP_206_199 & nP_198_191;
  assign nG_205_190 = nG_205_198 | (nP_205_198 & nG_197_190);
  assign nP_205_190 = nP_205_198 & nP_197_190;
  assign nG_204_189 = nG_204_197 | (nP_204_197 & nG_196_189);
  assign nP_204_189 = nP_204_197 & nP_196_189;
  assign nG_203_188 = nG_203_196 | (nP_203_196 & nG_195_188);
  assign nP_203_188 = nP_203_196 & nP_195_188;
  assign nG_202_187 = nG_202_195 | (nP_202_195 & nG_194_187);
  assign nP_202_187 = nP_202_195 & nP_194_187;
  assign nG_201_186 = nG_201_194 | (nP_201_194 & nG_193_186);
  assign nP_201_186 = nP_201_194 & nP_193_186;
  assign nG_200_185 = nG_200_193 | (nP_200_193 & nG_192_185);
  assign nP_200_185 = nP_200_193 & nP_192_185;
  assign nG_199_184 = nG_199_192 | (nP_199_192 & nG_191_184);
  assign nP_199_184 = nP_199_192 & nP_191_184;
  assign nG_198_183 = nG_198_191 | (nP_198_191 & nG_190_183);
  assign nP_198_183 = nP_198_191 & nP_190_183;
  assign nG_197_182 = nG_197_190 | (nP_197_190 & nG_189_182);
  assign nP_197_182 = nP_197_190 & nP_189_182;
  assign nG_196_181 = nG_196_189 | (nP_196_189 & nG_188_181);
  assign nP_196_181 = nP_196_189 & nP_188_181;
  assign nG_195_180 = nG_195_188 | (nP_195_188 & nG_187_180);
  assign nP_195_180 = nP_195_188 & nP_187_180;
  assign nG_194_179 = nG_194_187 | (nP_194_187 & nG_186_179);
  assign nP_194_179 = nP_194_187 & nP_186_179;
  assign nG_193_178 = nG_193_186 | (nP_193_186 & nG_185_178);
  assign nP_193_178 = nP_193_186 & nP_185_178;
  assign nG_192_177 = nG_192_185 | (nP_192_185 & nG_184_177);
  assign nP_192_177 = nP_192_185 & nP_184_177;
  assign nG_191_176 = nG_191_184 | (nP_191_184 & nG_183_176);
  assign nP_191_176 = nP_191_184 & nP_183_176;
  assign nG_190_175 = nG_190_183 | (nP_190_183 & nG_182_175);
  assign nP_190_175 = nP_190_183 & nP_182_175;
  assign nG_189_174 = nG_189_182 | (nP_189_182 & nG_181_174);
  assign nP_189_174 = nP_189_182 & nP_181_174;
  assign nG_188_173 = nG_188_181 | (nP_188_181 & nG_180_173);
  assign nP_188_173 = nP_188_181 & nP_180_173;
  assign nG_187_172 = nG_187_180 | (nP_187_180 & nG_179_172);
  assign nP_187_172 = nP_187_180 & nP_179_172;
  assign nG_186_171 = nG_186_179 | (nP_186_179 & nG_178_171);
  assign nP_186_171 = nP_186_179 & nP_178_171;
  assign nG_185_170 = nG_185_178 | (nP_185_178 & nG_177_170);
  assign nP_185_170 = nP_185_178 & nP_177_170;
  assign nG_184_169 = nG_184_177 | (nP_184_177 & nG_176_169);
  assign nP_184_169 = nP_184_177 & nP_176_169;
  assign nG_183_168 = nG_183_176 | (nP_183_176 & nG_175_168);
  assign nP_183_168 = nP_183_176 & nP_175_168;
  assign nG_182_167 = nG_182_175 | (nP_182_175 & nG_174_167);
  assign nP_182_167 = nP_182_175 & nP_174_167;
  assign nG_181_166 = nG_181_174 | (nP_181_174 & nG_173_166);
  assign nP_181_166 = nP_181_174 & nP_173_166;
  assign nG_180_165 = nG_180_173 | (nP_180_173 & nG_172_165);
  assign nP_180_165 = nP_180_173 & nP_172_165;
  assign nG_179_164 = nG_179_172 | (nP_179_172 & nG_171_164);
  assign nP_179_164 = nP_179_172 & nP_171_164;
  assign nG_178_163 = nG_178_171 | (nP_178_171 & nG_170_163);
  assign nP_178_163 = nP_178_171 & nP_170_163;
  assign nG_177_162 = nG_177_170 | (nP_177_170 & nG_169_162);
  assign nP_177_162 = nP_177_170 & nP_169_162;
  assign nG_176_161 = nG_176_169 | (nP_176_169 & nG_168_161);
  assign nP_176_161 = nP_176_169 & nP_168_161;
  assign nG_175_160 = nG_175_168 | (nP_175_168 & nG_167_160);
  assign nP_175_160 = nP_175_168 & nP_167_160;
  assign nG_174_159 = nG_174_167 | (nP_174_167 & nG_166_159);
  assign nP_174_159 = nP_174_167 & nP_166_159;
  assign nG_173_158 = nG_173_166 | (nP_173_166 & nG_165_158);
  assign nP_173_158 = nP_173_166 & nP_165_158;
  assign nG_172_157 = nG_172_165 | (nP_172_165 & nG_164_157);
  assign nP_172_157 = nP_172_165 & nP_164_157;
  assign nG_171_156 = nG_171_164 | (nP_171_164 & nG_163_156);
  assign nP_171_156 = nP_171_164 & nP_163_156;
  assign nG_170_155 = nG_170_163 | (nP_170_163 & nG_162_155);
  assign nP_170_155 = nP_170_163 & nP_162_155;
  assign nG_169_154 = nG_169_162 | (nP_169_162 & nG_161_154);
  assign nP_169_154 = nP_169_162 & nP_161_154;
  assign nG_168_153 = nG_168_161 | (nP_168_161 & nG_160_153);
  assign nP_168_153 = nP_168_161 & nP_160_153;
  assign nG_167_152 = nG_167_160 | (nP_167_160 & nG_159_152);
  assign nP_167_152 = nP_167_160 & nP_159_152;
  assign nG_166_151 = nG_166_159 | (nP_166_159 & nG_158_151);
  assign nP_166_151 = nP_166_159 & nP_158_151;
  assign nG_165_150 = nG_165_158 | (nP_165_158 & nG_157_150);
  assign nP_165_150 = nP_165_158 & nP_157_150;
  assign nG_164_149 = nG_164_157 | (nP_164_157 & nG_156_149);
  assign nP_164_149 = nP_164_157 & nP_156_149;
  assign nG_163_148 = nG_163_156 | (nP_163_156 & nG_155_148);
  assign nP_163_148 = nP_163_156 & nP_155_148;
  assign nG_162_147 = nG_162_155 | (nP_162_155 & nG_154_147);
  assign nP_162_147 = nP_162_155 & nP_154_147;
  assign nG_161_146 = nG_161_154 | (nP_161_154 & nG_153_146);
  assign nP_161_146 = nP_161_154 & nP_153_146;
  assign nG_160_145 = nG_160_153 | (nP_160_153 & nG_152_145);
  assign nP_160_145 = nP_160_153 & nP_152_145;
  assign nG_159_144 = nG_159_152 | (nP_159_152 & nG_151_144);
  assign nP_159_144 = nP_159_152 & nP_151_144;
  assign nG_158_143 = nG_158_151 | (nP_158_151 & nG_150_143);
  assign nP_158_143 = nP_158_151 & nP_150_143;
  assign nG_157_142 = nG_157_150 | (nP_157_150 & nG_149_142);
  assign nP_157_142 = nP_157_150 & nP_149_142;
  assign nG_156_141 = nG_156_149 | (nP_156_149 & nG_148_141);
  assign nP_156_141 = nP_156_149 & nP_148_141;
  assign nG_155_140 = nG_155_148 | (nP_155_148 & nG_147_140);
  assign nP_155_140 = nP_155_148 & nP_147_140;
  assign nG_154_139 = nG_154_147 | (nP_154_147 & nG_146_139);
  assign nP_154_139 = nP_154_147 & nP_146_139;
  assign nG_153_138 = nG_153_146 | (nP_153_146 & nG_145_138);
  assign nP_153_138 = nP_153_146 & nP_145_138;
  assign nG_152_137 = nG_152_145 | (nP_152_145 & nG_144_137);
  assign nP_152_137 = nP_152_145 & nP_144_137;
  assign nG_151_136 = nG_151_144 | (nP_151_144 & nG_143_136);
  assign nP_151_136 = nP_151_144 & nP_143_136;
  assign nG_150_135 = nG_150_143 | (nP_150_143 & nG_142_135);
  assign nP_150_135 = nP_150_143 & nP_142_135;
  assign nG_149_134 = nG_149_142 | (nP_149_142 & nG_141_134);
  assign nP_149_134 = nP_149_142 & nP_141_134;
  assign nG_148_133 = nG_148_141 | (nP_148_141 & nG_140_133);
  assign nP_148_133 = nP_148_141 & nP_140_133;
  assign nG_147_132 = nG_147_140 | (nP_147_140 & nG_139_132);
  assign nP_147_132 = nP_147_140 & nP_139_132;
  assign nG_146_131 = nG_146_139 | (nP_146_139 & nG_138_131);
  assign nP_146_131 = nP_146_139 & nP_138_131;
  assign nG_145_130 = nG_145_138 | (nP_145_138 & nG_137_130);
  assign nP_145_130 = nP_145_138 & nP_137_130;
  assign nG_144_129 = nG_144_137 | (nP_144_137 & nG_136_129);
  assign nP_144_129 = nP_144_137 & nP_136_129;
  assign nG_143_128 = nG_143_136 | (nP_143_136 & nG_135_128);
  assign nP_143_128 = nP_143_136 & nP_135_128;
  assign nG_142_127 = nG_142_135 | (nP_142_135 & nG_134_127);
  assign nP_142_127 = nP_142_135 & nP_134_127;
  assign nG_141_126 = nG_141_134 | (nP_141_134 & nG_133_126);
  assign nP_141_126 = nP_141_134 & nP_133_126;
  assign nG_140_125 = nG_140_133 | (nP_140_133 & nG_132_125);
  assign nP_140_125 = nP_140_133 & nP_132_125;
  assign nG_139_124 = nG_139_132 | (nP_139_132 & nG_131_124);
  assign nP_139_124 = nP_139_132 & nP_131_124;
  assign nG_138_123 = nG_138_131 | (nP_138_131 & nG_130_123);
  assign nP_138_123 = nP_138_131 & nP_130_123;
  assign nG_137_122 = nG_137_130 | (nP_137_130 & nG_129_122);
  assign nP_137_122 = nP_137_130 & nP_129_122;
  assign nG_136_121 = nG_136_129 | (nP_136_129 & nG_128_121);
  assign nP_136_121 = nP_136_129 & nP_128_121;
  assign nG_135_120 = nG_135_128 | (nP_135_128 & nG_127_120);
  assign nP_135_120 = nP_135_128 & nP_127_120;
  assign nG_134_119 = nG_134_127 | (nP_134_127 & nG_126_119);
  assign nP_134_119 = nP_134_127 & nP_126_119;
  assign nG_133_118 = nG_133_126 | (nP_133_126 & nG_125_118);
  assign nP_133_118 = nP_133_126 & nP_125_118;
  assign nG_132_117 = nG_132_125 | (nP_132_125 & nG_124_117);
  assign nP_132_117 = nP_132_125 & nP_124_117;
  assign nG_131_116 = nG_131_124 | (nP_131_124 & nG_123_116);
  assign nP_131_116 = nP_131_124 & nP_123_116;
  assign nG_130_115 = nG_130_123 | (nP_130_123 & nG_122_115);
  assign nP_130_115 = nP_130_123 & nP_122_115;
  assign nG_129_114 = nG_129_122 | (nP_129_122 & nG_121_114);
  assign nP_129_114 = nP_129_122 & nP_121_114;
  assign nG_128_113 = nG_128_121 | (nP_128_121 & nG_120_113);
  assign nP_128_113 = nP_128_121 & nP_120_113;
  assign nG_127_112 = nG_127_120 | (nP_127_120 & nG_119_112);
  assign nP_127_112 = nP_127_120 & nP_119_112;
  assign nG_126_111 = nG_126_119 | (nP_126_119 & nG_118_111);
  assign nP_126_111 = nP_126_119 & nP_118_111;
  assign nG_125_110 = nG_125_118 | (nP_125_118 & nG_117_110);
  assign nP_125_110 = nP_125_118 & nP_117_110;
  assign nG_124_109 = nG_124_117 | (nP_124_117 & nG_116_109);
  assign nP_124_109 = nP_124_117 & nP_116_109;
  assign nG_123_108 = nG_123_116 | (nP_123_116 & nG_115_108);
  assign nP_123_108 = nP_123_116 & nP_115_108;
  assign nG_122_107 = nG_122_115 | (nP_122_115 & nG_114_107);
  assign nP_122_107 = nP_122_115 & nP_114_107;
  assign nG_121_106 = nG_121_114 | (nP_121_114 & nG_113_106);
  assign nP_121_106 = nP_121_114 & nP_113_106;
  assign nG_120_105 = nG_120_113 | (nP_120_113 & nG_112_105);
  assign nP_120_105 = nP_120_113 & nP_112_105;
  assign nG_119_104 = nG_119_112 | (nP_119_112 & nG_111_104);
  assign nP_119_104 = nP_119_112 & nP_111_104;
  assign nG_118_103 = nG_118_111 | (nP_118_111 & nG_110_103);
  assign nP_118_103 = nP_118_111 & nP_110_103;
  assign nG_117_102 = nG_117_110 | (nP_117_110 & nG_109_102);
  assign nP_117_102 = nP_117_110 & nP_109_102;
  assign nG_116_101 = nG_116_109 | (nP_116_109 & nG_108_101);
  assign nP_116_101 = nP_116_109 & nP_108_101;
  assign nG_115_100 = nG_115_108 | (nP_115_108 & nG_107_100);
  assign nP_115_100 = nP_115_108 & nP_107_100;
  assign nG_114_99 = nG_114_107 | (nP_114_107 & nG_106_99);
  assign nP_114_99 = nP_114_107 & nP_106_99;
  assign nG_113_98 = nG_113_106 | (nP_113_106 & nG_105_98);
  assign nP_113_98 = nP_113_106 & nP_105_98;
  assign nG_112_97 = nG_112_105 | (nP_112_105 & nG_104_97);
  assign nP_112_97 = nP_112_105 & nP_104_97;
  assign nG_111_96 = nG_111_104 | (nP_111_104 & nG_103_96);
  assign nP_111_96 = nP_111_104 & nP_103_96;
  assign nG_110_95 = nG_110_103 | (nP_110_103 & nG_102_95);
  assign nP_110_95 = nP_110_103 & nP_102_95;
  assign nG_109_94 = nG_109_102 | (nP_109_102 & nG_101_94);
  assign nP_109_94 = nP_109_102 & nP_101_94;
  assign nG_108_93 = nG_108_101 | (nP_108_101 & nG_100_93);
  assign nP_108_93 = nP_108_101 & nP_100_93;
  assign nG_107_92 = nG_107_100 | (nP_107_100 & nG_99_92);
  assign nP_107_92 = nP_107_100 & nP_99_92;
  assign nG_106_91 = nG_106_99 | (nP_106_99 & nG_98_91);
  assign nP_106_91 = nP_106_99 & nP_98_91;
  assign nG_105_90 = nG_105_98 | (nP_105_98 & nG_97_90);
  assign nP_105_90 = nP_105_98 & nP_97_90;
  assign nG_104_89 = nG_104_97 | (nP_104_97 & nG_96_89);
  assign nP_104_89 = nP_104_97 & nP_96_89;
  assign nG_103_88 = nG_103_96 | (nP_103_96 & nG_95_88);
  assign nP_103_88 = nP_103_96 & nP_95_88;
  assign nG_102_87 = nG_102_95 | (nP_102_95 & nG_94_87);
  assign nP_102_87 = nP_102_95 & nP_94_87;
  assign nG_101_86 = nG_101_94 | (nP_101_94 & nG_93_86);
  assign nP_101_86 = nP_101_94 & nP_93_86;
  assign nG_100_85 = nG_100_93 | (nP_100_93 & nG_92_85);
  assign nP_100_85 = nP_100_93 & nP_92_85;
  assign nG_99_84 = nG_99_92 | (nP_99_92 & nG_91_84);
  assign nP_99_84 = nP_99_92 & nP_91_84;
  assign nG_98_83 = nG_98_91 | (nP_98_91 & nG_90_83);
  assign nP_98_83 = nP_98_91 & nP_90_83;
  assign nG_97_82 = nG_97_90 | (nP_97_90 & nG_89_82);
  assign nP_97_82 = nP_97_90 & nP_89_82;
  assign nG_96_81 = nG_96_89 | (nP_96_89 & nG_88_81);
  assign nP_96_81 = nP_96_89 & nP_88_81;
  assign nG_95_80 = nG_95_88 | (nP_95_88 & nG_87_80);
  assign nP_95_80 = nP_95_88 & nP_87_80;
  assign nG_94_79 = nG_94_87 | (nP_94_87 & nG_86_79);
  assign nP_94_79 = nP_94_87 & nP_86_79;
  assign nG_93_78 = nG_93_86 | (nP_93_86 & nG_85_78);
  assign nP_93_78 = nP_93_86 & nP_85_78;
  assign nG_92_77 = nG_92_85 | (nP_92_85 & nG_84_77);
  assign nP_92_77 = nP_92_85 & nP_84_77;
  assign nG_91_76 = nG_91_84 | (nP_91_84 & nG_83_76);
  assign nP_91_76 = nP_91_84 & nP_83_76;
  assign nG_90_75 = nG_90_83 | (nP_90_83 & nG_82_75);
  assign nP_90_75 = nP_90_83 & nP_82_75;
  assign nG_89_74 = nG_89_82 | (nP_89_82 & nG_81_74);
  assign nP_89_74 = nP_89_82 & nP_81_74;
  assign nG_88_73 = nG_88_81 | (nP_88_81 & nG_80_73);
  assign nP_88_73 = nP_88_81 & nP_80_73;
  assign nG_87_72 = nG_87_80 | (nP_87_80 & nG_79_72);
  assign nP_87_72 = nP_87_80 & nP_79_72;
  assign nG_86_71 = nG_86_79 | (nP_86_79 & nG_78_71);
  assign nP_86_71 = nP_86_79 & nP_78_71;
  assign nG_85_70 = nG_85_78 | (nP_85_78 & nG_77_70);
  assign nP_85_70 = nP_85_78 & nP_77_70;
  assign nG_84_69 = nG_84_77 | (nP_84_77 & nG_76_69);
  assign nP_84_69 = nP_84_77 & nP_76_69;
  assign nG_83_68 = nG_83_76 | (nP_83_76 & nG_75_68);
  assign nP_83_68 = nP_83_76 & nP_75_68;
  assign nG_82_67 = nG_82_75 | (nP_82_75 & nG_74_67);
  assign nP_82_67 = nP_82_75 & nP_74_67;
  assign nG_81_66 = nG_81_74 | (nP_81_74 & nG_73_66);
  assign nP_81_66 = nP_81_74 & nP_73_66;
  assign nG_80_65 = nG_80_73 | (nP_80_73 & nG_72_65);
  assign nP_80_65 = nP_80_73 & nP_72_65;
  assign nG_79_64 = nG_79_72 | (nP_79_72 & nG_71_64);
  assign nP_79_64 = nP_79_72 & nP_71_64;
  assign nG_78_63 = nG_78_71 | (nP_78_71 & nG_70_63);
  assign nP_78_63 = nP_78_71 & nP_70_63;
  assign nG_77_62 = nG_77_70 | (nP_77_70 & nG_69_62);
  assign nP_77_62 = nP_77_70 & nP_69_62;
  assign nG_76_61 = nG_76_69 | (nP_76_69 & nG_68_61);
  assign nP_76_61 = nP_76_69 & nP_68_61;
  assign nG_75_60 = nG_75_68 | (nP_75_68 & nG_67_60);
  assign nP_75_60 = nP_75_68 & nP_67_60;
  assign nG_74_59 = nG_74_67 | (nP_74_67 & nG_66_59);
  assign nP_74_59 = nP_74_67 & nP_66_59;
  assign nG_73_58 = nG_73_66 | (nP_73_66 & nG_65_58);
  assign nP_73_58 = nP_73_66 & nP_65_58;
  assign nG_72_57 = nG_72_65 | (nP_72_65 & nG_64_57);
  assign nP_72_57 = nP_72_65 & nP_64_57;
  assign nG_71_56 = nG_71_64 | (nP_71_64 & nG_63_56);
  assign nP_71_56 = nP_71_64 & nP_63_56;
  assign nG_70_55 = nG_70_63 | (nP_70_63 & nG_62_55);
  assign nP_70_55 = nP_70_63 & nP_62_55;
  assign nG_69_54 = nG_69_62 | (nP_69_62 & nG_61_54);
  assign nP_69_54 = nP_69_62 & nP_61_54;
  assign nG_68_53 = nG_68_61 | (nP_68_61 & nG_60_53);
  assign nP_68_53 = nP_68_61 & nP_60_53;
  assign nG_67_52 = nG_67_60 | (nP_67_60 & nG_59_52);
  assign nP_67_52 = nP_67_60 & nP_59_52;
  assign nG_66_51 = nG_66_59 | (nP_66_59 & nG_58_51);
  assign nP_66_51 = nP_66_59 & nP_58_51;
  assign nG_65_50 = nG_65_58 | (nP_65_58 & nG_57_50);
  assign nP_65_50 = nP_65_58 & nP_57_50;
  assign nG_64_49 = nG_64_57 | (nP_64_57 & nG_56_49);
  assign nP_64_49 = nP_64_57 & nP_56_49;
  assign nG_63_48 = nG_63_56 | (nP_63_56 & nG_55_48);
  assign nP_63_48 = nP_63_56 & nP_55_48;
  assign nG_62_47 = nG_62_55 | (nP_62_55 & nG_54_47);
  assign nP_62_47 = nP_62_55 & nP_54_47;
  assign nG_61_46 = nG_61_54 | (nP_61_54 & nG_53_46);
  assign nP_61_46 = nP_61_54 & nP_53_46;
  assign nG_60_45 = nG_60_53 | (nP_60_53 & nG_52_45);
  assign nP_60_45 = nP_60_53 & nP_52_45;
  assign nG_59_44 = nG_59_52 | (nP_59_52 & nG_51_44);
  assign nP_59_44 = nP_59_52 & nP_51_44;
  assign nG_58_43 = nG_58_51 | (nP_58_51 & nG_50_43);
  assign nP_58_43 = nP_58_51 & nP_50_43;
  assign nG_57_42 = nG_57_50 | (nP_57_50 & nG_49_42);
  assign nP_57_42 = nP_57_50 & nP_49_42;
  assign nG_56_41 = nG_56_49 | (nP_56_49 & nG_48_41);
  assign nP_56_41 = nP_56_49 & nP_48_41;
  assign nG_55_40 = nG_55_48 | (nP_55_48 & nG_47_40);
  assign nP_55_40 = nP_55_48 & nP_47_40;
  assign nG_54_39 = nG_54_47 | (nP_54_47 & nG_46_39);
  assign nP_54_39 = nP_54_47 & nP_46_39;
  assign nG_53_38 = nG_53_46 | (nP_53_46 & nG_45_38);
  assign nP_53_38 = nP_53_46 & nP_45_38;
  assign nG_52_37 = nG_52_45 | (nP_52_45 & nG_44_37);
  assign nP_52_37 = nP_52_45 & nP_44_37;
  assign nG_51_36 = nG_51_44 | (nP_51_44 & nG_43_36);
  assign nP_51_36 = nP_51_44 & nP_43_36;
  assign nG_50_35 = nG_50_43 | (nP_50_43 & nG_42_35);
  assign nP_50_35 = nP_50_43 & nP_42_35;
  assign nG_49_34 = nG_49_42 | (nP_49_42 & nG_41_34);
  assign nP_49_34 = nP_49_42 & nP_41_34;
  assign nG_48_33 = nG_48_41 | (nP_48_41 & nG_40_33);
  assign nP_48_33 = nP_48_41 & nP_40_33;
  assign nG_47_32 = nG_47_40 | (nP_47_40 & nG_39_32);
  assign nP_47_32 = nP_47_40 & nP_39_32;
  assign nG_46_31 = nG_46_39 | (nP_46_39 & nG_38_31);
  assign nP_46_31 = nP_46_39 & nP_38_31;
  assign nG_45_30 = nG_45_38 | (nP_45_38 & nG_37_30);
  assign nP_45_30 = nP_45_38 & nP_37_30;
  assign nG_44_29 = nG_44_37 | (nP_44_37 & nG_36_29);
  assign nP_44_29 = nP_44_37 & nP_36_29;
  assign nG_43_28 = nG_43_36 | (nP_43_36 & nG_35_28);
  assign nP_43_28 = nP_43_36 & nP_35_28;
  assign nG_42_27 = nG_42_35 | (nP_42_35 & nG_34_27);
  assign nP_42_27 = nP_42_35 & nP_34_27;
  assign nG_41_26 = nG_41_34 | (nP_41_34 & nG_33_26);
  assign nP_41_26 = nP_41_34 & nP_33_26;
  assign nG_40_25 = nG_40_33 | (nP_40_33 & nG_32_25);
  assign nP_40_25 = nP_40_33 & nP_32_25;
  assign nG_39_24 = nG_39_32 | (nP_39_32 & nG_31_24);
  assign nP_39_24 = nP_39_32 & nP_31_24;
  assign nG_38_23 = nG_38_31 | (nP_38_31 & nG_30_23);
  assign nP_38_23 = nP_38_31 & nP_30_23;
  assign nG_37_22 = nG_37_30 | (nP_37_30 & nG_29_22);
  assign nP_37_22 = nP_37_30 & nP_29_22;
  assign nG_36_21 = nG_36_29 | (nP_36_29 & nG_28_21);
  assign nP_36_21 = nP_36_29 & nP_28_21;
  assign nG_35_20 = nG_35_28 | (nP_35_28 & nG_27_20);
  assign nP_35_20 = nP_35_28 & nP_27_20;
  assign nG_34_19 = nG_34_27 | (nP_34_27 & nG_26_19);
  assign nP_34_19 = nP_34_27 & nP_26_19;
  assign nG_33_18 = nG_33_26 | (nP_33_26 & nG_25_18);
  assign nP_33_18 = nP_33_26 & nP_25_18;
  assign nG_32_17 = nG_32_25 | (nP_32_25 & nG_24_17);
  assign nP_32_17 = nP_32_25 & nP_24_17;
  assign nG_31_16 = nG_31_24 | (nP_31_24 & nG_23_16);
  assign nP_31_16 = nP_31_24 & nP_23_16;
  assign nG_30_15 = nG_30_23 | (nP_30_23 & nG_22_15);
  assign nP_30_15 = nP_30_23 & nP_22_15;
  assign nG_29_14 = nG_29_22 | (nP_29_22 & nG_21_14);
  assign nP_29_14 = nP_29_22 & nP_21_14;
  assign nG_28_13 = nG_28_21 | (nP_28_21 & nG_20_13);
  assign nP_28_13 = nP_28_21 & nP_20_13;
  assign nG_27_12 = nG_27_20 | (nP_27_20 & nG_19_12);
  assign nP_27_12 = nP_27_20 & nP_19_12;
  assign nG_26_11 = nG_26_19 | (nP_26_19 & nG_18_11);
  assign nP_26_11 = nP_26_19 & nP_18_11;
  assign nG_25_10 = nG_25_18 | (nP_25_18 & nG_17_10);
  assign nP_25_10 = nP_25_18 & nP_17_10;
  assign nG_24_9 = nG_24_17 | (nP_24_17 & nG_16_9);
  assign nP_24_9 = nP_24_17 & nP_16_9;
  assign nG_23_8 = nG_23_16 | (nP_23_16 & nG_15_8);
  assign nP_23_8 = nP_23_16 & nP_15_8;
  assign nG_22_7 = nG_22_15 | (nP_22_15 & nG_14_7);
  assign nP_22_7 = nP_22_15 & nP_14_7;
  assign nG_21_6 = nG_21_14 | (nP_21_14 & nG_13_6);
  assign nP_21_6 = nP_21_14 & nP_13_6;
  assign nG_20_5 = nG_20_13 | (nP_20_13 & nG_12_5);
  assign nP_20_5 = nP_20_13 & nP_12_5;
  assign nG_19_4 = nG_19_12 | (nP_19_12 & nG_11_4);
  assign nP_19_4 = nP_19_12 & nP_11_4;
  assign nG_18_3 = nG_18_11 | (nP_18_11 & nG_10_3);
  assign nP_18_3 = nP_18_11 & nP_10_3;
  assign nG_17_2 = nG_17_10 | (nP_17_10 & nG_9_2);
  assign nP_17_2 = nP_17_10 & nP_9_2;
  assign nG_16_1 = nG_16_9 | (nP_16_9 & nG_8_1);
  assign nP_16_1 = nP_16_9 & nP_8_1;
  assign nG_15_0 = nG_15_8 | (nP_15_8 & nG_7_0);
  assign nP_15_0 = nP_15_8 & nP_7_0;
  assign nG_14_0 = nG_14_7 | (nP_14_7 & nG_6_0);
  assign nP_14_0 = nP_14_7 & nP_6_0;
  assign nG_13_0 = nG_13_6 | (nP_13_6 & nG_5_0);
  assign nP_13_0 = nP_13_6 & nP_5_0;
  assign nG_12_0 = nG_12_5 | (nP_12_5 & nG_4_0);
  assign nP_12_0 = nP_12_5 & nP_4_0;
  assign nG_11_0 = nG_11_4 | (nP_11_4 & nG_3_0);
  assign nP_11_0 = nP_11_4 & nP_3_0;
  assign nG_10_0 = nG_10_3 | (nP_10_3 & nG_2_0);
  assign nP_10_0 = nP_10_3 & nP_2_0;
  assign nG_9_0 = nG_9_2 | (nP_9_2 & nG_1_0);
  assign nP_9_0 = nP_9_2 & nP_1_0;
  assign nG_8_0 = nG_8_1 | (nP_8_1 & nG_0_0);
  assign nP_8_0 = nP_8_1 & nP_0_0;

  assign nG_255_224 = nG_255_240 | (nP_255_240 & nG_239_224);
  assign nP_255_224 = nP_255_240 & nP_239_224;
  assign nG_254_223 = nG_254_239 | (nP_254_239 & nG_238_223);
  assign nP_254_223 = nP_254_239 & nP_238_223;
  assign nG_253_222 = nG_253_238 | (nP_253_238 & nG_237_222);
  assign nP_253_222 = nP_253_238 & nP_237_222;
  assign nG_252_221 = nG_252_237 | (nP_252_237 & nG_236_221);
  assign nP_252_221 = nP_252_237 & nP_236_221;
  assign nG_251_220 = nG_251_236 | (nP_251_236 & nG_235_220);
  assign nP_251_220 = nP_251_236 & nP_235_220;
  assign nG_250_219 = nG_250_235 | (nP_250_235 & nG_234_219);
  assign nP_250_219 = nP_250_235 & nP_234_219;
  assign nG_249_218 = nG_249_234 | (nP_249_234 & nG_233_218);
  assign nP_249_218 = nP_249_234 & nP_233_218;
  assign nG_248_217 = nG_248_233 | (nP_248_233 & nG_232_217);
  assign nP_248_217 = nP_248_233 & nP_232_217;
  assign nG_247_216 = nG_247_232 | (nP_247_232 & nG_231_216);
  assign nP_247_216 = nP_247_232 & nP_231_216;
  assign nG_246_215 = nG_246_231 | (nP_246_231 & nG_230_215);
  assign nP_246_215 = nP_246_231 & nP_230_215;
  assign nG_245_214 = nG_245_230 | (nP_245_230 & nG_229_214);
  assign nP_245_214 = nP_245_230 & nP_229_214;
  assign nG_244_213 = nG_244_229 | (nP_244_229 & nG_228_213);
  assign nP_244_213 = nP_244_229 & nP_228_213;
  assign nG_243_212 = nG_243_228 | (nP_243_228 & nG_227_212);
  assign nP_243_212 = nP_243_228 & nP_227_212;
  assign nG_242_211 = nG_242_227 | (nP_242_227 & nG_226_211);
  assign nP_242_211 = nP_242_227 & nP_226_211;
  assign nG_241_210 = nG_241_226 | (nP_241_226 & nG_225_210);
  assign nP_241_210 = nP_241_226 & nP_225_210;
  assign nG_240_209 = nG_240_225 | (nP_240_225 & nG_224_209);
  assign nP_240_209 = nP_240_225 & nP_224_209;
  assign nG_239_208 = nG_239_224 | (nP_239_224 & nG_223_208);
  assign nP_239_208 = nP_239_224 & nP_223_208;
  assign nG_238_207 = nG_238_223 | (nP_238_223 & nG_222_207);
  assign nP_238_207 = nP_238_223 & nP_222_207;
  assign nG_237_206 = nG_237_222 | (nP_237_222 & nG_221_206);
  assign nP_237_206 = nP_237_222 & nP_221_206;
  assign nG_236_205 = nG_236_221 | (nP_236_221 & nG_220_205);
  assign nP_236_205 = nP_236_221 & nP_220_205;
  assign nG_235_204 = nG_235_220 | (nP_235_220 & nG_219_204);
  assign nP_235_204 = nP_235_220 & nP_219_204;
  assign nG_234_203 = nG_234_219 | (nP_234_219 & nG_218_203);
  assign nP_234_203 = nP_234_219 & nP_218_203;
  assign nG_233_202 = nG_233_218 | (nP_233_218 & nG_217_202);
  assign nP_233_202 = nP_233_218 & nP_217_202;
  assign nG_232_201 = nG_232_217 | (nP_232_217 & nG_216_201);
  assign nP_232_201 = nP_232_217 & nP_216_201;
  assign nG_231_200 = nG_231_216 | (nP_231_216 & nG_215_200);
  assign nP_231_200 = nP_231_216 & nP_215_200;
  assign nG_230_199 = nG_230_215 | (nP_230_215 & nG_214_199);
  assign nP_230_199 = nP_230_215 & nP_214_199;
  assign nG_229_198 = nG_229_214 | (nP_229_214 & nG_213_198);
  assign nP_229_198 = nP_229_214 & nP_213_198;
  assign nG_228_197 = nG_228_213 | (nP_228_213 & nG_212_197);
  assign nP_228_197 = nP_228_213 & nP_212_197;
  assign nG_227_196 = nG_227_212 | (nP_227_212 & nG_211_196);
  assign nP_227_196 = nP_227_212 & nP_211_196;
  assign nG_226_195 = nG_226_211 | (nP_226_211 & nG_210_195);
  assign nP_226_195 = nP_226_211 & nP_210_195;
  assign nG_225_194 = nG_225_210 | (nP_225_210 & nG_209_194);
  assign nP_225_194 = nP_225_210 & nP_209_194;
  assign nG_224_193 = nG_224_209 | (nP_224_209 & nG_208_193);
  assign nP_224_193 = nP_224_209 & nP_208_193;
  assign nG_223_192 = nG_223_208 | (nP_223_208 & nG_207_192);
  assign nP_223_192 = nP_223_208 & nP_207_192;
  assign nG_222_191 = nG_222_207 | (nP_222_207 & nG_206_191);
  assign nP_222_191 = nP_222_207 & nP_206_191;
  assign nG_221_190 = nG_221_206 | (nP_221_206 & nG_205_190);
  assign nP_221_190 = nP_221_206 & nP_205_190;
  assign nG_220_189 = nG_220_205 | (nP_220_205 & nG_204_189);
  assign nP_220_189 = nP_220_205 & nP_204_189;
  assign nG_219_188 = nG_219_204 | (nP_219_204 & nG_203_188);
  assign nP_219_188 = nP_219_204 & nP_203_188;
  assign nG_218_187 = nG_218_203 | (nP_218_203 & nG_202_187);
  assign nP_218_187 = nP_218_203 & nP_202_187;
  assign nG_217_186 = nG_217_202 | (nP_217_202 & nG_201_186);
  assign nP_217_186 = nP_217_202 & nP_201_186;
  assign nG_216_185 = nG_216_201 | (nP_216_201 & nG_200_185);
  assign nP_216_185 = nP_216_201 & nP_200_185;
  assign nG_215_184 = nG_215_200 | (nP_215_200 & nG_199_184);
  assign nP_215_184 = nP_215_200 & nP_199_184;
  assign nG_214_183 = nG_214_199 | (nP_214_199 & nG_198_183);
  assign nP_214_183 = nP_214_199 & nP_198_183;
  assign nG_213_182 = nG_213_198 | (nP_213_198 & nG_197_182);
  assign nP_213_182 = nP_213_198 & nP_197_182;
  assign nG_212_181 = nG_212_197 | (nP_212_197 & nG_196_181);
  assign nP_212_181 = nP_212_197 & nP_196_181;
  assign nG_211_180 = nG_211_196 | (nP_211_196 & nG_195_180);
  assign nP_211_180 = nP_211_196 & nP_195_180;
  assign nG_210_179 = nG_210_195 | (nP_210_195 & nG_194_179);
  assign nP_210_179 = nP_210_195 & nP_194_179;
  assign nG_209_178 = nG_209_194 | (nP_209_194 & nG_193_178);
  assign nP_209_178 = nP_209_194 & nP_193_178;
  assign nG_208_177 = nG_208_193 | (nP_208_193 & nG_192_177);
  assign nP_208_177 = nP_208_193 & nP_192_177;
  assign nG_207_176 = nG_207_192 | (nP_207_192 & nG_191_176);
  assign nP_207_176 = nP_207_192 & nP_191_176;
  assign nG_206_175 = nG_206_191 | (nP_206_191 & nG_190_175);
  assign nP_206_175 = nP_206_191 & nP_190_175;
  assign nG_205_174 = nG_205_190 | (nP_205_190 & nG_189_174);
  assign nP_205_174 = nP_205_190 & nP_189_174;
  assign nG_204_173 = nG_204_189 | (nP_204_189 & nG_188_173);
  assign nP_204_173 = nP_204_189 & nP_188_173;
  assign nG_203_172 = nG_203_188 | (nP_203_188 & nG_187_172);
  assign nP_203_172 = nP_203_188 & nP_187_172;
  assign nG_202_171 = nG_202_187 | (nP_202_187 & nG_186_171);
  assign nP_202_171 = nP_202_187 & nP_186_171;
  assign nG_201_170 = nG_201_186 | (nP_201_186 & nG_185_170);
  assign nP_201_170 = nP_201_186 & nP_185_170;
  assign nG_200_169 = nG_200_185 | (nP_200_185 & nG_184_169);
  assign nP_200_169 = nP_200_185 & nP_184_169;
  assign nG_199_168 = nG_199_184 | (nP_199_184 & nG_183_168);
  assign nP_199_168 = nP_199_184 & nP_183_168;
  assign nG_198_167 = nG_198_183 | (nP_198_183 & nG_182_167);
  assign nP_198_167 = nP_198_183 & nP_182_167;
  assign nG_197_166 = nG_197_182 | (nP_197_182 & nG_181_166);
  assign nP_197_166 = nP_197_182 & nP_181_166;
  assign nG_196_165 = nG_196_181 | (nP_196_181 & nG_180_165);
  assign nP_196_165 = nP_196_181 & nP_180_165;
  assign nG_195_164 = nG_195_180 | (nP_195_180 & nG_179_164);
  assign nP_195_164 = nP_195_180 & nP_179_164;
  assign nG_194_163 = nG_194_179 | (nP_194_179 & nG_178_163);
  assign nP_194_163 = nP_194_179 & nP_178_163;
  assign nG_193_162 = nG_193_178 | (nP_193_178 & nG_177_162);
  assign nP_193_162 = nP_193_178 & nP_177_162;
  assign nG_192_161 = nG_192_177 | (nP_192_177 & nG_176_161);
  assign nP_192_161 = nP_192_177 & nP_176_161;
  assign nG_191_160 = nG_191_176 | (nP_191_176 & nG_175_160);
  assign nP_191_160 = nP_191_176 & nP_175_160;
  assign nG_190_159 = nG_190_175 | (nP_190_175 & nG_174_159);
  assign nP_190_159 = nP_190_175 & nP_174_159;
  assign nG_189_158 = nG_189_174 | (nP_189_174 & nG_173_158);
  assign nP_189_158 = nP_189_174 & nP_173_158;
  assign nG_188_157 = nG_188_173 | (nP_188_173 & nG_172_157);
  assign nP_188_157 = nP_188_173 & nP_172_157;
  assign nG_187_156 = nG_187_172 | (nP_187_172 & nG_171_156);
  assign nP_187_156 = nP_187_172 & nP_171_156;
  assign nG_186_155 = nG_186_171 | (nP_186_171 & nG_170_155);
  assign nP_186_155 = nP_186_171 & nP_170_155;
  assign nG_185_154 = nG_185_170 | (nP_185_170 & nG_169_154);
  assign nP_185_154 = nP_185_170 & nP_169_154;
  assign nG_184_153 = nG_184_169 | (nP_184_169 & nG_168_153);
  assign nP_184_153 = nP_184_169 & nP_168_153;
  assign nG_183_152 = nG_183_168 | (nP_183_168 & nG_167_152);
  assign nP_183_152 = nP_183_168 & nP_167_152;
  assign nG_182_151 = nG_182_167 | (nP_182_167 & nG_166_151);
  assign nP_182_151 = nP_182_167 & nP_166_151;
  assign nG_181_150 = nG_181_166 | (nP_181_166 & nG_165_150);
  assign nP_181_150 = nP_181_166 & nP_165_150;
  assign nG_180_149 = nG_180_165 | (nP_180_165 & nG_164_149);
  assign nP_180_149 = nP_180_165 & nP_164_149;
  assign nG_179_148 = nG_179_164 | (nP_179_164 & nG_163_148);
  assign nP_179_148 = nP_179_164 & nP_163_148;
  assign nG_178_147 = nG_178_163 | (nP_178_163 & nG_162_147);
  assign nP_178_147 = nP_178_163 & nP_162_147;
  assign nG_177_146 = nG_177_162 | (nP_177_162 & nG_161_146);
  assign nP_177_146 = nP_177_162 & nP_161_146;
  assign nG_176_145 = nG_176_161 | (nP_176_161 & nG_160_145);
  assign nP_176_145 = nP_176_161 & nP_160_145;
  assign nG_175_144 = nG_175_160 | (nP_175_160 & nG_159_144);
  assign nP_175_144 = nP_175_160 & nP_159_144;
  assign nG_174_143 = nG_174_159 | (nP_174_159 & nG_158_143);
  assign nP_174_143 = nP_174_159 & nP_158_143;
  assign nG_173_142 = nG_173_158 | (nP_173_158 & nG_157_142);
  assign nP_173_142 = nP_173_158 & nP_157_142;
  assign nG_172_141 = nG_172_157 | (nP_172_157 & nG_156_141);
  assign nP_172_141 = nP_172_157 & nP_156_141;
  assign nG_171_140 = nG_171_156 | (nP_171_156 & nG_155_140);
  assign nP_171_140 = nP_171_156 & nP_155_140;
  assign nG_170_139 = nG_170_155 | (nP_170_155 & nG_154_139);
  assign nP_170_139 = nP_170_155 & nP_154_139;
  assign nG_169_138 = nG_169_154 | (nP_169_154 & nG_153_138);
  assign nP_169_138 = nP_169_154 & nP_153_138;
  assign nG_168_137 = nG_168_153 | (nP_168_153 & nG_152_137);
  assign nP_168_137 = nP_168_153 & nP_152_137;
  assign nG_167_136 = nG_167_152 | (nP_167_152 & nG_151_136);
  assign nP_167_136 = nP_167_152 & nP_151_136;
  assign nG_166_135 = nG_166_151 | (nP_166_151 & nG_150_135);
  assign nP_166_135 = nP_166_151 & nP_150_135;
  assign nG_165_134 = nG_165_150 | (nP_165_150 & nG_149_134);
  assign nP_165_134 = nP_165_150 & nP_149_134;
  assign nG_164_133 = nG_164_149 | (nP_164_149 & nG_148_133);
  assign nP_164_133 = nP_164_149 & nP_148_133;
  assign nG_163_132 = nG_163_148 | (nP_163_148 & nG_147_132);
  assign nP_163_132 = nP_163_148 & nP_147_132;
  assign nG_162_131 = nG_162_147 | (nP_162_147 & nG_146_131);
  assign nP_162_131 = nP_162_147 & nP_146_131;
  assign nG_161_130 = nG_161_146 | (nP_161_146 & nG_145_130);
  assign nP_161_130 = nP_161_146 & nP_145_130;
  assign nG_160_129 = nG_160_145 | (nP_160_145 & nG_144_129);
  assign nP_160_129 = nP_160_145 & nP_144_129;
  assign nG_159_128 = nG_159_144 | (nP_159_144 & nG_143_128);
  assign nP_159_128 = nP_159_144 & nP_143_128;
  assign nG_158_127 = nG_158_143 | (nP_158_143 & nG_142_127);
  assign nP_158_127 = nP_158_143 & nP_142_127;
  assign nG_157_126 = nG_157_142 | (nP_157_142 & nG_141_126);
  assign nP_157_126 = nP_157_142 & nP_141_126;
  assign nG_156_125 = nG_156_141 | (nP_156_141 & nG_140_125);
  assign nP_156_125 = nP_156_141 & nP_140_125;
  assign nG_155_124 = nG_155_140 | (nP_155_140 & nG_139_124);
  assign nP_155_124 = nP_155_140 & nP_139_124;
  assign nG_154_123 = nG_154_139 | (nP_154_139 & nG_138_123);
  assign nP_154_123 = nP_154_139 & nP_138_123;
  assign nG_153_122 = nG_153_138 | (nP_153_138 & nG_137_122);
  assign nP_153_122 = nP_153_138 & nP_137_122;
  assign nG_152_121 = nG_152_137 | (nP_152_137 & nG_136_121);
  assign nP_152_121 = nP_152_137 & nP_136_121;
  assign nG_151_120 = nG_151_136 | (nP_151_136 & nG_135_120);
  assign nP_151_120 = nP_151_136 & nP_135_120;
  assign nG_150_119 = nG_150_135 | (nP_150_135 & nG_134_119);
  assign nP_150_119 = nP_150_135 & nP_134_119;
  assign nG_149_118 = nG_149_134 | (nP_149_134 & nG_133_118);
  assign nP_149_118 = nP_149_134 & nP_133_118;
  assign nG_148_117 = nG_148_133 | (nP_148_133 & nG_132_117);
  assign nP_148_117 = nP_148_133 & nP_132_117;
  assign nG_147_116 = nG_147_132 | (nP_147_132 & nG_131_116);
  assign nP_147_116 = nP_147_132 & nP_131_116;
  assign nG_146_115 = nG_146_131 | (nP_146_131 & nG_130_115);
  assign nP_146_115 = nP_146_131 & nP_130_115;
  assign nG_145_114 = nG_145_130 | (nP_145_130 & nG_129_114);
  assign nP_145_114 = nP_145_130 & nP_129_114;
  assign nG_144_113 = nG_144_129 | (nP_144_129 & nG_128_113);
  assign nP_144_113 = nP_144_129 & nP_128_113;
  assign nG_143_112 = nG_143_128 | (nP_143_128 & nG_127_112);
  assign nP_143_112 = nP_143_128 & nP_127_112;
  assign nG_142_111 = nG_142_127 | (nP_142_127 & nG_126_111);
  assign nP_142_111 = nP_142_127 & nP_126_111;
  assign nG_141_110 = nG_141_126 | (nP_141_126 & nG_125_110);
  assign nP_141_110 = nP_141_126 & nP_125_110;
  assign nG_140_109 = nG_140_125 | (nP_140_125 & nG_124_109);
  assign nP_140_109 = nP_140_125 & nP_124_109;
  assign nG_139_108 = nG_139_124 | (nP_139_124 & nG_123_108);
  assign nP_139_108 = nP_139_124 & nP_123_108;
  assign nG_138_107 = nG_138_123 | (nP_138_123 & nG_122_107);
  assign nP_138_107 = nP_138_123 & nP_122_107;
  assign nG_137_106 = nG_137_122 | (nP_137_122 & nG_121_106);
  assign nP_137_106 = nP_137_122 & nP_121_106;
  assign nG_136_105 = nG_136_121 | (nP_136_121 & nG_120_105);
  assign nP_136_105 = nP_136_121 & nP_120_105;
  assign nG_135_104 = nG_135_120 | (nP_135_120 & nG_119_104);
  assign nP_135_104 = nP_135_120 & nP_119_104;
  assign nG_134_103 = nG_134_119 | (nP_134_119 & nG_118_103);
  assign nP_134_103 = nP_134_119 & nP_118_103;
  assign nG_133_102 = nG_133_118 | (nP_133_118 & nG_117_102);
  assign nP_133_102 = nP_133_118 & nP_117_102;
  assign nG_132_101 = nG_132_117 | (nP_132_117 & nG_116_101);
  assign nP_132_101 = nP_132_117 & nP_116_101;
  assign nG_131_100 = nG_131_116 | (nP_131_116 & nG_115_100);
  assign nP_131_100 = nP_131_116 & nP_115_100;
  assign nG_130_99 = nG_130_115 | (nP_130_115 & nG_114_99);
  assign nP_130_99 = nP_130_115 & nP_114_99;
  assign nG_129_98 = nG_129_114 | (nP_129_114 & nG_113_98);
  assign nP_129_98 = nP_129_114 & nP_113_98;
  assign nG_128_97 = nG_128_113 | (nP_128_113 & nG_112_97);
  assign nP_128_97 = nP_128_113 & nP_112_97;
  assign nG_127_96 = nG_127_112 | (nP_127_112 & nG_111_96);
  assign nP_127_96 = nP_127_112 & nP_111_96;
  assign nG_126_95 = nG_126_111 | (nP_126_111 & nG_110_95);
  assign nP_126_95 = nP_126_111 & nP_110_95;
  assign nG_125_94 = nG_125_110 | (nP_125_110 & nG_109_94);
  assign nP_125_94 = nP_125_110 & nP_109_94;
  assign nG_124_93 = nG_124_109 | (nP_124_109 & nG_108_93);
  assign nP_124_93 = nP_124_109 & nP_108_93;
  assign nG_123_92 = nG_123_108 | (nP_123_108 & nG_107_92);
  assign nP_123_92 = nP_123_108 & nP_107_92;
  assign nG_122_91 = nG_122_107 | (nP_122_107 & nG_106_91);
  assign nP_122_91 = nP_122_107 & nP_106_91;
  assign nG_121_90 = nG_121_106 | (nP_121_106 & nG_105_90);
  assign nP_121_90 = nP_121_106 & nP_105_90;
  assign nG_120_89 = nG_120_105 | (nP_120_105 & nG_104_89);
  assign nP_120_89 = nP_120_105 & nP_104_89;
  assign nG_119_88 = nG_119_104 | (nP_119_104 & nG_103_88);
  assign nP_119_88 = nP_119_104 & nP_103_88;
  assign nG_118_87 = nG_118_103 | (nP_118_103 & nG_102_87);
  assign nP_118_87 = nP_118_103 & nP_102_87;
  assign nG_117_86 = nG_117_102 | (nP_117_102 & nG_101_86);
  assign nP_117_86 = nP_117_102 & nP_101_86;
  assign nG_116_85 = nG_116_101 | (nP_116_101 & nG_100_85);
  assign nP_116_85 = nP_116_101 & nP_100_85;
  assign nG_115_84 = nG_115_100 | (nP_115_100 & nG_99_84);
  assign nP_115_84 = nP_115_100 & nP_99_84;
  assign nG_114_83 = nG_114_99 | (nP_114_99 & nG_98_83);
  assign nP_114_83 = nP_114_99 & nP_98_83;
  assign nG_113_82 = nG_113_98 | (nP_113_98 & nG_97_82);
  assign nP_113_82 = nP_113_98 & nP_97_82;
  assign nG_112_81 = nG_112_97 | (nP_112_97 & nG_96_81);
  assign nP_112_81 = nP_112_97 & nP_96_81;
  assign nG_111_80 = nG_111_96 | (nP_111_96 & nG_95_80);
  assign nP_111_80 = nP_111_96 & nP_95_80;
  assign nG_110_79 = nG_110_95 | (nP_110_95 & nG_94_79);
  assign nP_110_79 = nP_110_95 & nP_94_79;
  assign nG_109_78 = nG_109_94 | (nP_109_94 & nG_93_78);
  assign nP_109_78 = nP_109_94 & nP_93_78;
  assign nG_108_77 = nG_108_93 | (nP_108_93 & nG_92_77);
  assign nP_108_77 = nP_108_93 & nP_92_77;
  assign nG_107_76 = nG_107_92 | (nP_107_92 & nG_91_76);
  assign nP_107_76 = nP_107_92 & nP_91_76;
  assign nG_106_75 = nG_106_91 | (nP_106_91 & nG_90_75);
  assign nP_106_75 = nP_106_91 & nP_90_75;
  assign nG_105_74 = nG_105_90 | (nP_105_90 & nG_89_74);
  assign nP_105_74 = nP_105_90 & nP_89_74;
  assign nG_104_73 = nG_104_89 | (nP_104_89 & nG_88_73);
  assign nP_104_73 = nP_104_89 & nP_88_73;
  assign nG_103_72 = nG_103_88 | (nP_103_88 & nG_87_72);
  assign nP_103_72 = nP_103_88 & nP_87_72;
  assign nG_102_71 = nG_102_87 | (nP_102_87 & nG_86_71);
  assign nP_102_71 = nP_102_87 & nP_86_71;
  assign nG_101_70 = nG_101_86 | (nP_101_86 & nG_85_70);
  assign nP_101_70 = nP_101_86 & nP_85_70;
  assign nG_100_69 = nG_100_85 | (nP_100_85 & nG_84_69);
  assign nP_100_69 = nP_100_85 & nP_84_69;
  assign nG_99_68 = nG_99_84 | (nP_99_84 & nG_83_68);
  assign nP_99_68 = nP_99_84 & nP_83_68;
  assign nG_98_67 = nG_98_83 | (nP_98_83 & nG_82_67);
  assign nP_98_67 = nP_98_83 & nP_82_67;
  assign nG_97_66 = nG_97_82 | (nP_97_82 & nG_81_66);
  assign nP_97_66 = nP_97_82 & nP_81_66;
  assign nG_96_65 = nG_96_81 | (nP_96_81 & nG_80_65);
  assign nP_96_65 = nP_96_81 & nP_80_65;
  assign nG_95_64 = nG_95_80 | (nP_95_80 & nG_79_64);
  assign nP_95_64 = nP_95_80 & nP_79_64;
  assign nG_94_63 = nG_94_79 | (nP_94_79 & nG_78_63);
  assign nP_94_63 = nP_94_79 & nP_78_63;
  assign nG_93_62 = nG_93_78 | (nP_93_78 & nG_77_62);
  assign nP_93_62 = nP_93_78 & nP_77_62;
  assign nG_92_61 = nG_92_77 | (nP_92_77 & nG_76_61);
  assign nP_92_61 = nP_92_77 & nP_76_61;
  assign nG_91_60 = nG_91_76 | (nP_91_76 & nG_75_60);
  assign nP_91_60 = nP_91_76 & nP_75_60;
  assign nG_90_59 = nG_90_75 | (nP_90_75 & nG_74_59);
  assign nP_90_59 = nP_90_75 & nP_74_59;
  assign nG_89_58 = nG_89_74 | (nP_89_74 & nG_73_58);
  assign nP_89_58 = nP_89_74 & nP_73_58;
  assign nG_88_57 = nG_88_73 | (nP_88_73 & nG_72_57);
  assign nP_88_57 = nP_88_73 & nP_72_57;
  assign nG_87_56 = nG_87_72 | (nP_87_72 & nG_71_56);
  assign nP_87_56 = nP_87_72 & nP_71_56;
  assign nG_86_55 = nG_86_71 | (nP_86_71 & nG_70_55);
  assign nP_86_55 = nP_86_71 & nP_70_55;
  assign nG_85_54 = nG_85_70 | (nP_85_70 & nG_69_54);
  assign nP_85_54 = nP_85_70 & nP_69_54;
  assign nG_84_53 = nG_84_69 | (nP_84_69 & nG_68_53);
  assign nP_84_53 = nP_84_69 & nP_68_53;
  assign nG_83_52 = nG_83_68 | (nP_83_68 & nG_67_52);
  assign nP_83_52 = nP_83_68 & nP_67_52;
  assign nG_82_51 = nG_82_67 | (nP_82_67 & nG_66_51);
  assign nP_82_51 = nP_82_67 & nP_66_51;
  assign nG_81_50 = nG_81_66 | (nP_81_66 & nG_65_50);
  assign nP_81_50 = nP_81_66 & nP_65_50;
  assign nG_80_49 = nG_80_65 | (nP_80_65 & nG_64_49);
  assign nP_80_49 = nP_80_65 & nP_64_49;
  assign nG_79_48 = nG_79_64 | (nP_79_64 & nG_63_48);
  assign nP_79_48 = nP_79_64 & nP_63_48;
  assign nG_78_47 = nG_78_63 | (nP_78_63 & nG_62_47);
  assign nP_78_47 = nP_78_63 & nP_62_47;
  assign nG_77_46 = nG_77_62 | (nP_77_62 & nG_61_46);
  assign nP_77_46 = nP_77_62 & nP_61_46;
  assign nG_76_45 = nG_76_61 | (nP_76_61 & nG_60_45);
  assign nP_76_45 = nP_76_61 & nP_60_45;
  assign nG_75_44 = nG_75_60 | (nP_75_60 & nG_59_44);
  assign nP_75_44 = nP_75_60 & nP_59_44;
  assign nG_74_43 = nG_74_59 | (nP_74_59 & nG_58_43);
  assign nP_74_43 = nP_74_59 & nP_58_43;
  assign nG_73_42 = nG_73_58 | (nP_73_58 & nG_57_42);
  assign nP_73_42 = nP_73_58 & nP_57_42;
  assign nG_72_41 = nG_72_57 | (nP_72_57 & nG_56_41);
  assign nP_72_41 = nP_72_57 & nP_56_41;
  assign nG_71_40 = nG_71_56 | (nP_71_56 & nG_55_40);
  assign nP_71_40 = nP_71_56 & nP_55_40;
  assign nG_70_39 = nG_70_55 | (nP_70_55 & nG_54_39);
  assign nP_70_39 = nP_70_55 & nP_54_39;
  assign nG_69_38 = nG_69_54 | (nP_69_54 & nG_53_38);
  assign nP_69_38 = nP_69_54 & nP_53_38;
  assign nG_68_37 = nG_68_53 | (nP_68_53 & nG_52_37);
  assign nP_68_37 = nP_68_53 & nP_52_37;
  assign nG_67_36 = nG_67_52 | (nP_67_52 & nG_51_36);
  assign nP_67_36 = nP_67_52 & nP_51_36;
  assign nG_66_35 = nG_66_51 | (nP_66_51 & nG_50_35);
  assign nP_66_35 = nP_66_51 & nP_50_35;
  assign nG_65_34 = nG_65_50 | (nP_65_50 & nG_49_34);
  assign nP_65_34 = nP_65_50 & nP_49_34;
  assign nG_64_33 = nG_64_49 | (nP_64_49 & nG_48_33);
  assign nP_64_33 = nP_64_49 & nP_48_33;
  assign nG_63_32 = nG_63_48 | (nP_63_48 & nG_47_32);
  assign nP_63_32 = nP_63_48 & nP_47_32;
  assign nG_62_31 = nG_62_47 | (nP_62_47 & nG_46_31);
  assign nP_62_31 = nP_62_47 & nP_46_31;
  assign nG_61_30 = nG_61_46 | (nP_61_46 & nG_45_30);
  assign nP_61_30 = nP_61_46 & nP_45_30;
  assign nG_60_29 = nG_60_45 | (nP_60_45 & nG_44_29);
  assign nP_60_29 = nP_60_45 & nP_44_29;
  assign nG_59_28 = nG_59_44 | (nP_59_44 & nG_43_28);
  assign nP_59_28 = nP_59_44 & nP_43_28;
  assign nG_58_27 = nG_58_43 | (nP_58_43 & nG_42_27);
  assign nP_58_27 = nP_58_43 & nP_42_27;
  assign nG_57_26 = nG_57_42 | (nP_57_42 & nG_41_26);
  assign nP_57_26 = nP_57_42 & nP_41_26;
  assign nG_56_25 = nG_56_41 | (nP_56_41 & nG_40_25);
  assign nP_56_25 = nP_56_41 & nP_40_25;
  assign nG_55_24 = nG_55_40 | (nP_55_40 & nG_39_24);
  assign nP_55_24 = nP_55_40 & nP_39_24;
  assign nG_54_23 = nG_54_39 | (nP_54_39 & nG_38_23);
  assign nP_54_23 = nP_54_39 & nP_38_23;
  assign nG_53_22 = nG_53_38 | (nP_53_38 & nG_37_22);
  assign nP_53_22 = nP_53_38 & nP_37_22;
  assign nG_52_21 = nG_52_37 | (nP_52_37 & nG_36_21);
  assign nP_52_21 = nP_52_37 & nP_36_21;
  assign nG_51_20 = nG_51_36 | (nP_51_36 & nG_35_20);
  assign nP_51_20 = nP_51_36 & nP_35_20;
  assign nG_50_19 = nG_50_35 | (nP_50_35 & nG_34_19);
  assign nP_50_19 = nP_50_35 & nP_34_19;
  assign nG_49_18 = nG_49_34 | (nP_49_34 & nG_33_18);
  assign nP_49_18 = nP_49_34 & nP_33_18;
  assign nG_48_17 = nG_48_33 | (nP_48_33 & nG_32_17);
  assign nP_48_17 = nP_48_33 & nP_32_17;
  assign nG_47_16 = nG_47_32 | (nP_47_32 & nG_31_16);
  assign nP_47_16 = nP_47_32 & nP_31_16;
  assign nG_46_15 = nG_46_31 | (nP_46_31 & nG_30_15);
  assign nP_46_15 = nP_46_31 & nP_30_15;
  assign nG_45_14 = nG_45_30 | (nP_45_30 & nG_29_14);
  assign nP_45_14 = nP_45_30 & nP_29_14;
  assign nG_44_13 = nG_44_29 | (nP_44_29 & nG_28_13);
  assign nP_44_13 = nP_44_29 & nP_28_13;
  assign nG_43_12 = nG_43_28 | (nP_43_28 & nG_27_12);
  assign nP_43_12 = nP_43_28 & nP_27_12;
  assign nG_42_11 = nG_42_27 | (nP_42_27 & nG_26_11);
  assign nP_42_11 = nP_42_27 & nP_26_11;
  assign nG_41_10 = nG_41_26 | (nP_41_26 & nG_25_10);
  assign nP_41_10 = nP_41_26 & nP_25_10;
  assign nG_40_9 = nG_40_25 | (nP_40_25 & nG_24_9);
  assign nP_40_9 = nP_40_25 & nP_24_9;
  assign nG_39_8 = nG_39_24 | (nP_39_24 & nG_23_8);
  assign nP_39_8 = nP_39_24 & nP_23_8;
  assign nG_38_7 = nG_38_23 | (nP_38_23 & nG_22_7);
  assign nP_38_7 = nP_38_23 & nP_22_7;
  assign nG_37_6 = nG_37_22 | (nP_37_22 & nG_21_6);
  assign nP_37_6 = nP_37_22 & nP_21_6;
  assign nG_36_5 = nG_36_21 | (nP_36_21 & nG_20_5);
  assign nP_36_5 = nP_36_21 & nP_20_5;
  assign nG_35_4 = nG_35_20 | (nP_35_20 & nG_19_4);
  assign nP_35_4 = nP_35_20 & nP_19_4;
  assign nG_34_3 = nG_34_19 | (nP_34_19 & nG_18_3);
  assign nP_34_3 = nP_34_19 & nP_18_3;
  assign nG_33_2 = nG_33_18 | (nP_33_18 & nG_17_2);
  assign nP_33_2 = nP_33_18 & nP_17_2;
  assign nG_32_1 = nG_32_17 | (nP_32_17 & nG_16_1);
  assign nP_32_1 = nP_32_17 & nP_16_1;
  assign nG_31_0 = nG_31_16 | (nP_31_16 & nG_15_0);
  assign nP_31_0 = nP_31_16 & nP_15_0;
  assign nG_30_0 = nG_30_15 | (nP_30_15 & nG_14_0);
  assign nP_30_0 = nP_30_15 & nP_14_0;
  assign nG_29_0 = nG_29_14 | (nP_29_14 & nG_13_0);
  assign nP_29_0 = nP_29_14 & nP_13_0;
  assign nG_28_0 = nG_28_13 | (nP_28_13 & nG_12_0);
  assign nP_28_0 = nP_28_13 & nP_12_0;
  assign nG_27_0 = nG_27_12 | (nP_27_12 & nG_11_0);
  assign nP_27_0 = nP_27_12 & nP_11_0;
  assign nG_26_0 = nG_26_11 | (nP_26_11 & nG_10_0);
  assign nP_26_0 = nP_26_11 & nP_10_0;
  assign nG_25_0 = nG_25_10 | (nP_25_10 & nG_9_0);
  assign nP_25_0 = nP_25_10 & nP_9_0;
  assign nG_24_0 = nG_24_9 | (nP_24_9 & nG_8_0);
  assign nP_24_0 = nP_24_9 & nP_8_0;
  assign nG_23_0 = nG_23_8 | (nP_23_8 & nG_7_0);
  assign nP_23_0 = nP_23_8 & nP_7_0;
  assign nG_22_0 = nG_22_7 | (nP_22_7 & nG_6_0);
  assign nP_22_0 = nP_22_7 & nP_6_0;
  assign nG_21_0 = nG_21_6 | (nP_21_6 & nG_5_0);
  assign nP_21_0 = nP_21_6 & nP_5_0;
  assign nG_20_0 = nG_20_5 | (nP_20_5 & nG_4_0);
  assign nP_20_0 = nP_20_5 & nP_4_0;
  assign nG_19_0 = nG_19_4 | (nP_19_4 & nG_3_0);
  assign nP_19_0 = nP_19_4 & nP_3_0;
  assign nG_18_0 = nG_18_3 | (nP_18_3 & nG_2_0);
  assign nP_18_0 = nP_18_3 & nP_2_0;
  assign nG_17_0 = nG_17_2 | (nP_17_2 & nG_1_0);
  assign nP_17_0 = nP_17_2 & nP_1_0;
  assign nG_16_0 = nG_16_1 | (nP_16_1 & nG_0_0);
  assign nP_16_0 = nP_16_1 & nP_0_0;

  assign nG_255_192 = nG_255_224 | (nP_255_224 & nG_223_192);
  assign nP_255_192 = nP_255_224 & nP_223_192;
  assign nG_254_191 = nG_254_223 | (nP_254_223 & nG_222_191);
  assign nP_254_191 = nP_254_223 & nP_222_191;
  assign nG_253_190 = nG_253_222 | (nP_253_222 & nG_221_190);
  assign nP_253_190 = nP_253_222 & nP_221_190;
  assign nG_252_189 = nG_252_221 | (nP_252_221 & nG_220_189);
  assign nP_252_189 = nP_252_221 & nP_220_189;
  assign nG_251_188 = nG_251_220 | (nP_251_220 & nG_219_188);
  assign nP_251_188 = nP_251_220 & nP_219_188;
  assign nG_250_187 = nG_250_219 | (nP_250_219 & nG_218_187);
  assign nP_250_187 = nP_250_219 & nP_218_187;
  assign nG_249_186 = nG_249_218 | (nP_249_218 & nG_217_186);
  assign nP_249_186 = nP_249_218 & nP_217_186;
  assign nG_248_185 = nG_248_217 | (nP_248_217 & nG_216_185);
  assign nP_248_185 = nP_248_217 & nP_216_185;
  assign nG_247_184 = nG_247_216 | (nP_247_216 & nG_215_184);
  assign nP_247_184 = nP_247_216 & nP_215_184;
  assign nG_246_183 = nG_246_215 | (nP_246_215 & nG_214_183);
  assign nP_246_183 = nP_246_215 & nP_214_183;
  assign nG_245_182 = nG_245_214 | (nP_245_214 & nG_213_182);
  assign nP_245_182 = nP_245_214 & nP_213_182;
  assign nG_244_181 = nG_244_213 | (nP_244_213 & nG_212_181);
  assign nP_244_181 = nP_244_213 & nP_212_181;
  assign nG_243_180 = nG_243_212 | (nP_243_212 & nG_211_180);
  assign nP_243_180 = nP_243_212 & nP_211_180;
  assign nG_242_179 = nG_242_211 | (nP_242_211 & nG_210_179);
  assign nP_242_179 = nP_242_211 & nP_210_179;
  assign nG_241_178 = nG_241_210 | (nP_241_210 & nG_209_178);
  assign nP_241_178 = nP_241_210 & nP_209_178;
  assign nG_240_177 = nG_240_209 | (nP_240_209 & nG_208_177);
  assign nP_240_177 = nP_240_209 & nP_208_177;
  assign nG_239_176 = nG_239_208 | (nP_239_208 & nG_207_176);
  assign nP_239_176 = nP_239_208 & nP_207_176;
  assign nG_238_175 = nG_238_207 | (nP_238_207 & nG_206_175);
  assign nP_238_175 = nP_238_207 & nP_206_175;
  assign nG_237_174 = nG_237_206 | (nP_237_206 & nG_205_174);
  assign nP_237_174 = nP_237_206 & nP_205_174;
  assign nG_236_173 = nG_236_205 | (nP_236_205 & nG_204_173);
  assign nP_236_173 = nP_236_205 & nP_204_173;
  assign nG_235_172 = nG_235_204 | (nP_235_204 & nG_203_172);
  assign nP_235_172 = nP_235_204 & nP_203_172;
  assign nG_234_171 = nG_234_203 | (nP_234_203 & nG_202_171);
  assign nP_234_171 = nP_234_203 & nP_202_171;
  assign nG_233_170 = nG_233_202 | (nP_233_202 & nG_201_170);
  assign nP_233_170 = nP_233_202 & nP_201_170;
  assign nG_232_169 = nG_232_201 | (nP_232_201 & nG_200_169);
  assign nP_232_169 = nP_232_201 & nP_200_169;
  assign nG_231_168 = nG_231_200 | (nP_231_200 & nG_199_168);
  assign nP_231_168 = nP_231_200 & nP_199_168;
  assign nG_230_167 = nG_230_199 | (nP_230_199 & nG_198_167);
  assign nP_230_167 = nP_230_199 & nP_198_167;
  assign nG_229_166 = nG_229_198 | (nP_229_198 & nG_197_166);
  assign nP_229_166 = nP_229_198 & nP_197_166;
  assign nG_228_165 = nG_228_197 | (nP_228_197 & nG_196_165);
  assign nP_228_165 = nP_228_197 & nP_196_165;
  assign nG_227_164 = nG_227_196 | (nP_227_196 & nG_195_164);
  assign nP_227_164 = nP_227_196 & nP_195_164;
  assign nG_226_163 = nG_226_195 | (nP_226_195 & nG_194_163);
  assign nP_226_163 = nP_226_195 & nP_194_163;
  assign nG_225_162 = nG_225_194 | (nP_225_194 & nG_193_162);
  assign nP_225_162 = nP_225_194 & nP_193_162;
  assign nG_224_161 = nG_224_193 | (nP_224_193 & nG_192_161);
  assign nP_224_161 = nP_224_193 & nP_192_161;
  assign nG_223_160 = nG_223_192 | (nP_223_192 & nG_191_160);
  assign nP_223_160 = nP_223_192 & nP_191_160;
  assign nG_222_159 = nG_222_191 | (nP_222_191 & nG_190_159);
  assign nP_222_159 = nP_222_191 & nP_190_159;
  assign nG_221_158 = nG_221_190 | (nP_221_190 & nG_189_158);
  assign nP_221_158 = nP_221_190 & nP_189_158;
  assign nG_220_157 = nG_220_189 | (nP_220_189 & nG_188_157);
  assign nP_220_157 = nP_220_189 & nP_188_157;
  assign nG_219_156 = nG_219_188 | (nP_219_188 & nG_187_156);
  assign nP_219_156 = nP_219_188 & nP_187_156;
  assign nG_218_155 = nG_218_187 | (nP_218_187 & nG_186_155);
  assign nP_218_155 = nP_218_187 & nP_186_155;
  assign nG_217_154 = nG_217_186 | (nP_217_186 & nG_185_154);
  assign nP_217_154 = nP_217_186 & nP_185_154;
  assign nG_216_153 = nG_216_185 | (nP_216_185 & nG_184_153);
  assign nP_216_153 = nP_216_185 & nP_184_153;
  assign nG_215_152 = nG_215_184 | (nP_215_184 & nG_183_152);
  assign nP_215_152 = nP_215_184 & nP_183_152;
  assign nG_214_151 = nG_214_183 | (nP_214_183 & nG_182_151);
  assign nP_214_151 = nP_214_183 & nP_182_151;
  assign nG_213_150 = nG_213_182 | (nP_213_182 & nG_181_150);
  assign nP_213_150 = nP_213_182 & nP_181_150;
  assign nG_212_149 = nG_212_181 | (nP_212_181 & nG_180_149);
  assign nP_212_149 = nP_212_181 & nP_180_149;
  assign nG_211_148 = nG_211_180 | (nP_211_180 & nG_179_148);
  assign nP_211_148 = nP_211_180 & nP_179_148;
  assign nG_210_147 = nG_210_179 | (nP_210_179 & nG_178_147);
  assign nP_210_147 = nP_210_179 & nP_178_147;
  assign nG_209_146 = nG_209_178 | (nP_209_178 & nG_177_146);
  assign nP_209_146 = nP_209_178 & nP_177_146;
  assign nG_208_145 = nG_208_177 | (nP_208_177 & nG_176_145);
  assign nP_208_145 = nP_208_177 & nP_176_145;
  assign nG_207_144 = nG_207_176 | (nP_207_176 & nG_175_144);
  assign nP_207_144 = nP_207_176 & nP_175_144;
  assign nG_206_143 = nG_206_175 | (nP_206_175 & nG_174_143);
  assign nP_206_143 = nP_206_175 & nP_174_143;
  assign nG_205_142 = nG_205_174 | (nP_205_174 & nG_173_142);
  assign nP_205_142 = nP_205_174 & nP_173_142;
  assign nG_204_141 = nG_204_173 | (nP_204_173 & nG_172_141);
  assign nP_204_141 = nP_204_173 & nP_172_141;
  assign nG_203_140 = nG_203_172 | (nP_203_172 & nG_171_140);
  assign nP_203_140 = nP_203_172 & nP_171_140;
  assign nG_202_139 = nG_202_171 | (nP_202_171 & nG_170_139);
  assign nP_202_139 = nP_202_171 & nP_170_139;
  assign nG_201_138 = nG_201_170 | (nP_201_170 & nG_169_138);
  assign nP_201_138 = nP_201_170 & nP_169_138;
  assign nG_200_137 = nG_200_169 | (nP_200_169 & nG_168_137);
  assign nP_200_137 = nP_200_169 & nP_168_137;
  assign nG_199_136 = nG_199_168 | (nP_199_168 & nG_167_136);
  assign nP_199_136 = nP_199_168 & nP_167_136;
  assign nG_198_135 = nG_198_167 | (nP_198_167 & nG_166_135);
  assign nP_198_135 = nP_198_167 & nP_166_135;
  assign nG_197_134 = nG_197_166 | (nP_197_166 & nG_165_134);
  assign nP_197_134 = nP_197_166 & nP_165_134;
  assign nG_196_133 = nG_196_165 | (nP_196_165 & nG_164_133);
  assign nP_196_133 = nP_196_165 & nP_164_133;
  assign nG_195_132 = nG_195_164 | (nP_195_164 & nG_163_132);
  assign nP_195_132 = nP_195_164 & nP_163_132;
  assign nG_194_131 = nG_194_163 | (nP_194_163 & nG_162_131);
  assign nP_194_131 = nP_194_163 & nP_162_131;
  assign nG_193_130 = nG_193_162 | (nP_193_162 & nG_161_130);
  assign nP_193_130 = nP_193_162 & nP_161_130;
  assign nG_192_129 = nG_192_161 | (nP_192_161 & nG_160_129);
  assign nP_192_129 = nP_192_161 & nP_160_129;
  assign nG_191_128 = nG_191_160 | (nP_191_160 & nG_159_128);
  assign nP_191_128 = nP_191_160 & nP_159_128;
  assign nG_190_127 = nG_190_159 | (nP_190_159 & nG_158_127);
  assign nP_190_127 = nP_190_159 & nP_158_127;
  assign nG_189_126 = nG_189_158 | (nP_189_158 & nG_157_126);
  assign nP_189_126 = nP_189_158 & nP_157_126;
  assign nG_188_125 = nG_188_157 | (nP_188_157 & nG_156_125);
  assign nP_188_125 = nP_188_157 & nP_156_125;
  assign nG_187_124 = nG_187_156 | (nP_187_156 & nG_155_124);
  assign nP_187_124 = nP_187_156 & nP_155_124;
  assign nG_186_123 = nG_186_155 | (nP_186_155 & nG_154_123);
  assign nP_186_123 = nP_186_155 & nP_154_123;
  assign nG_185_122 = nG_185_154 | (nP_185_154 & nG_153_122);
  assign nP_185_122 = nP_185_154 & nP_153_122;
  assign nG_184_121 = nG_184_153 | (nP_184_153 & nG_152_121);
  assign nP_184_121 = nP_184_153 & nP_152_121;
  assign nG_183_120 = nG_183_152 | (nP_183_152 & nG_151_120);
  assign nP_183_120 = nP_183_152 & nP_151_120;
  assign nG_182_119 = nG_182_151 | (nP_182_151 & nG_150_119);
  assign nP_182_119 = nP_182_151 & nP_150_119;
  assign nG_181_118 = nG_181_150 | (nP_181_150 & nG_149_118);
  assign nP_181_118 = nP_181_150 & nP_149_118;
  assign nG_180_117 = nG_180_149 | (nP_180_149 & nG_148_117);
  assign nP_180_117 = nP_180_149 & nP_148_117;
  assign nG_179_116 = nG_179_148 | (nP_179_148 & nG_147_116);
  assign nP_179_116 = nP_179_148 & nP_147_116;
  assign nG_178_115 = nG_178_147 | (nP_178_147 & nG_146_115);
  assign nP_178_115 = nP_178_147 & nP_146_115;
  assign nG_177_114 = nG_177_146 | (nP_177_146 & nG_145_114);
  assign nP_177_114 = nP_177_146 & nP_145_114;
  assign nG_176_113 = nG_176_145 | (nP_176_145 & nG_144_113);
  assign nP_176_113 = nP_176_145 & nP_144_113;
  assign nG_175_112 = nG_175_144 | (nP_175_144 & nG_143_112);
  assign nP_175_112 = nP_175_144 & nP_143_112;
  assign nG_174_111 = nG_174_143 | (nP_174_143 & nG_142_111);
  assign nP_174_111 = nP_174_143 & nP_142_111;
  assign nG_173_110 = nG_173_142 | (nP_173_142 & nG_141_110);
  assign nP_173_110 = nP_173_142 & nP_141_110;
  assign nG_172_109 = nG_172_141 | (nP_172_141 & nG_140_109);
  assign nP_172_109 = nP_172_141 & nP_140_109;
  assign nG_171_108 = nG_171_140 | (nP_171_140 & nG_139_108);
  assign nP_171_108 = nP_171_140 & nP_139_108;
  assign nG_170_107 = nG_170_139 | (nP_170_139 & nG_138_107);
  assign nP_170_107 = nP_170_139 & nP_138_107;
  assign nG_169_106 = nG_169_138 | (nP_169_138 & nG_137_106);
  assign nP_169_106 = nP_169_138 & nP_137_106;
  assign nG_168_105 = nG_168_137 | (nP_168_137 & nG_136_105);
  assign nP_168_105 = nP_168_137 & nP_136_105;
  assign nG_167_104 = nG_167_136 | (nP_167_136 & nG_135_104);
  assign nP_167_104 = nP_167_136 & nP_135_104;
  assign nG_166_103 = nG_166_135 | (nP_166_135 & nG_134_103);
  assign nP_166_103 = nP_166_135 & nP_134_103;
  assign nG_165_102 = nG_165_134 | (nP_165_134 & nG_133_102);
  assign nP_165_102 = nP_165_134 & nP_133_102;
  assign nG_164_101 = nG_164_133 | (nP_164_133 & nG_132_101);
  assign nP_164_101 = nP_164_133 & nP_132_101;
  assign nG_163_100 = nG_163_132 | (nP_163_132 & nG_131_100);
  assign nP_163_100 = nP_163_132 & nP_131_100;
  assign nG_162_99 = nG_162_131 | (nP_162_131 & nG_130_99);
  assign nP_162_99 = nP_162_131 & nP_130_99;
  assign nG_161_98 = nG_161_130 | (nP_161_130 & nG_129_98);
  assign nP_161_98 = nP_161_130 & nP_129_98;
  assign nG_160_97 = nG_160_129 | (nP_160_129 & nG_128_97);
  assign nP_160_97 = nP_160_129 & nP_128_97;
  assign nG_159_96 = nG_159_128 | (nP_159_128 & nG_127_96);
  assign nP_159_96 = nP_159_128 & nP_127_96;
  assign nG_158_95 = nG_158_127 | (nP_158_127 & nG_126_95);
  assign nP_158_95 = nP_158_127 & nP_126_95;
  assign nG_157_94 = nG_157_126 | (nP_157_126 & nG_125_94);
  assign nP_157_94 = nP_157_126 & nP_125_94;
  assign nG_156_93 = nG_156_125 | (nP_156_125 & nG_124_93);
  assign nP_156_93 = nP_156_125 & nP_124_93;
  assign nG_155_92 = nG_155_124 | (nP_155_124 & nG_123_92);
  assign nP_155_92 = nP_155_124 & nP_123_92;
  assign nG_154_91 = nG_154_123 | (nP_154_123 & nG_122_91);
  assign nP_154_91 = nP_154_123 & nP_122_91;
  assign nG_153_90 = nG_153_122 | (nP_153_122 & nG_121_90);
  assign nP_153_90 = nP_153_122 & nP_121_90;
  assign nG_152_89 = nG_152_121 | (nP_152_121 & nG_120_89);
  assign nP_152_89 = nP_152_121 & nP_120_89;
  assign nG_151_88 = nG_151_120 | (nP_151_120 & nG_119_88);
  assign nP_151_88 = nP_151_120 & nP_119_88;
  assign nG_150_87 = nG_150_119 | (nP_150_119 & nG_118_87);
  assign nP_150_87 = nP_150_119 & nP_118_87;
  assign nG_149_86 = nG_149_118 | (nP_149_118 & nG_117_86);
  assign nP_149_86 = nP_149_118 & nP_117_86;
  assign nG_148_85 = nG_148_117 | (nP_148_117 & nG_116_85);
  assign nP_148_85 = nP_148_117 & nP_116_85;
  assign nG_147_84 = nG_147_116 | (nP_147_116 & nG_115_84);
  assign nP_147_84 = nP_147_116 & nP_115_84;
  assign nG_146_83 = nG_146_115 | (nP_146_115 & nG_114_83);
  assign nP_146_83 = nP_146_115 & nP_114_83;
  assign nG_145_82 = nG_145_114 | (nP_145_114 & nG_113_82);
  assign nP_145_82 = nP_145_114 & nP_113_82;
  assign nG_144_81 = nG_144_113 | (nP_144_113 & nG_112_81);
  assign nP_144_81 = nP_144_113 & nP_112_81;
  assign nG_143_80 = nG_143_112 | (nP_143_112 & nG_111_80);
  assign nP_143_80 = nP_143_112 & nP_111_80;
  assign nG_142_79 = nG_142_111 | (nP_142_111 & nG_110_79);
  assign nP_142_79 = nP_142_111 & nP_110_79;
  assign nG_141_78 = nG_141_110 | (nP_141_110 & nG_109_78);
  assign nP_141_78 = nP_141_110 & nP_109_78;
  assign nG_140_77 = nG_140_109 | (nP_140_109 & nG_108_77);
  assign nP_140_77 = nP_140_109 & nP_108_77;
  assign nG_139_76 = nG_139_108 | (nP_139_108 & nG_107_76);
  assign nP_139_76 = nP_139_108 & nP_107_76;
  assign nG_138_75 = nG_138_107 | (nP_138_107 & nG_106_75);
  assign nP_138_75 = nP_138_107 & nP_106_75;
  assign nG_137_74 = nG_137_106 | (nP_137_106 & nG_105_74);
  assign nP_137_74 = nP_137_106 & nP_105_74;
  assign nG_136_73 = nG_136_105 | (nP_136_105 & nG_104_73);
  assign nP_136_73 = nP_136_105 & nP_104_73;
  assign nG_135_72 = nG_135_104 | (nP_135_104 & nG_103_72);
  assign nP_135_72 = nP_135_104 & nP_103_72;
  assign nG_134_71 = nG_134_103 | (nP_134_103 & nG_102_71);
  assign nP_134_71 = nP_134_103 & nP_102_71;
  assign nG_133_70 = nG_133_102 | (nP_133_102 & nG_101_70);
  assign nP_133_70 = nP_133_102 & nP_101_70;
  assign nG_132_69 = nG_132_101 | (nP_132_101 & nG_100_69);
  assign nP_132_69 = nP_132_101 & nP_100_69;
  assign nG_131_68 = nG_131_100 | (nP_131_100 & nG_99_68);
  assign nP_131_68 = nP_131_100 & nP_99_68;
  assign nG_130_67 = nG_130_99 | (nP_130_99 & nG_98_67);
  assign nP_130_67 = nP_130_99 & nP_98_67;
  assign nG_129_66 = nG_129_98 | (nP_129_98 & nG_97_66);
  assign nP_129_66 = nP_129_98 & nP_97_66;
  assign nG_128_65 = nG_128_97 | (nP_128_97 & nG_96_65);
  assign nP_128_65 = nP_128_97 & nP_96_65;
  assign nG_127_64 = nG_127_96 | (nP_127_96 & nG_95_64);
  assign nP_127_64 = nP_127_96 & nP_95_64;
  assign nG_126_63 = nG_126_95 | (nP_126_95 & nG_94_63);
  assign nP_126_63 = nP_126_95 & nP_94_63;
  assign nG_125_62 = nG_125_94 | (nP_125_94 & nG_93_62);
  assign nP_125_62 = nP_125_94 & nP_93_62;
  assign nG_124_61 = nG_124_93 | (nP_124_93 & nG_92_61);
  assign nP_124_61 = nP_124_93 & nP_92_61;
  assign nG_123_60 = nG_123_92 | (nP_123_92 & nG_91_60);
  assign nP_123_60 = nP_123_92 & nP_91_60;
  assign nG_122_59 = nG_122_91 | (nP_122_91 & nG_90_59);
  assign nP_122_59 = nP_122_91 & nP_90_59;
  assign nG_121_58 = nG_121_90 | (nP_121_90 & nG_89_58);
  assign nP_121_58 = nP_121_90 & nP_89_58;
  assign nG_120_57 = nG_120_89 | (nP_120_89 & nG_88_57);
  assign nP_120_57 = nP_120_89 & nP_88_57;
  assign nG_119_56 = nG_119_88 | (nP_119_88 & nG_87_56);
  assign nP_119_56 = nP_119_88 & nP_87_56;
  assign nG_118_55 = nG_118_87 | (nP_118_87 & nG_86_55);
  assign nP_118_55 = nP_118_87 & nP_86_55;
  assign nG_117_54 = nG_117_86 | (nP_117_86 & nG_85_54);
  assign nP_117_54 = nP_117_86 & nP_85_54;
  assign nG_116_53 = nG_116_85 | (nP_116_85 & nG_84_53);
  assign nP_116_53 = nP_116_85 & nP_84_53;
  assign nG_115_52 = nG_115_84 | (nP_115_84 & nG_83_52);
  assign nP_115_52 = nP_115_84 & nP_83_52;
  assign nG_114_51 = nG_114_83 | (nP_114_83 & nG_82_51);
  assign nP_114_51 = nP_114_83 & nP_82_51;
  assign nG_113_50 = nG_113_82 | (nP_113_82 & nG_81_50);
  assign nP_113_50 = nP_113_82 & nP_81_50;
  assign nG_112_49 = nG_112_81 | (nP_112_81 & nG_80_49);
  assign nP_112_49 = nP_112_81 & nP_80_49;
  assign nG_111_48 = nG_111_80 | (nP_111_80 & nG_79_48);
  assign nP_111_48 = nP_111_80 & nP_79_48;
  assign nG_110_47 = nG_110_79 | (nP_110_79 & nG_78_47);
  assign nP_110_47 = nP_110_79 & nP_78_47;
  assign nG_109_46 = nG_109_78 | (nP_109_78 & nG_77_46);
  assign nP_109_46 = nP_109_78 & nP_77_46;
  assign nG_108_45 = nG_108_77 | (nP_108_77 & nG_76_45);
  assign nP_108_45 = nP_108_77 & nP_76_45;
  assign nG_107_44 = nG_107_76 | (nP_107_76 & nG_75_44);
  assign nP_107_44 = nP_107_76 & nP_75_44;
  assign nG_106_43 = nG_106_75 | (nP_106_75 & nG_74_43);
  assign nP_106_43 = nP_106_75 & nP_74_43;
  assign nG_105_42 = nG_105_74 | (nP_105_74 & nG_73_42);
  assign nP_105_42 = nP_105_74 & nP_73_42;
  assign nG_104_41 = nG_104_73 | (nP_104_73 & nG_72_41);
  assign nP_104_41 = nP_104_73 & nP_72_41;
  assign nG_103_40 = nG_103_72 | (nP_103_72 & nG_71_40);
  assign nP_103_40 = nP_103_72 & nP_71_40;
  assign nG_102_39 = nG_102_71 | (nP_102_71 & nG_70_39);
  assign nP_102_39 = nP_102_71 & nP_70_39;
  assign nG_101_38 = nG_101_70 | (nP_101_70 & nG_69_38);
  assign nP_101_38 = nP_101_70 & nP_69_38;
  assign nG_100_37 = nG_100_69 | (nP_100_69 & nG_68_37);
  assign nP_100_37 = nP_100_69 & nP_68_37;
  assign nG_99_36 = nG_99_68 | (nP_99_68 & nG_67_36);
  assign nP_99_36 = nP_99_68 & nP_67_36;
  assign nG_98_35 = nG_98_67 | (nP_98_67 & nG_66_35);
  assign nP_98_35 = nP_98_67 & nP_66_35;
  assign nG_97_34 = nG_97_66 | (nP_97_66 & nG_65_34);
  assign nP_97_34 = nP_97_66 & nP_65_34;
  assign nG_96_33 = nG_96_65 | (nP_96_65 & nG_64_33);
  assign nP_96_33 = nP_96_65 & nP_64_33;
  assign nG_95_32 = nG_95_64 | (nP_95_64 & nG_63_32);
  assign nP_95_32 = nP_95_64 & nP_63_32;
  assign nG_94_31 = nG_94_63 | (nP_94_63 & nG_62_31);
  assign nP_94_31 = nP_94_63 & nP_62_31;
  assign nG_93_30 = nG_93_62 | (nP_93_62 & nG_61_30);
  assign nP_93_30 = nP_93_62 & nP_61_30;
  assign nG_92_29 = nG_92_61 | (nP_92_61 & nG_60_29);
  assign nP_92_29 = nP_92_61 & nP_60_29;
  assign nG_91_28 = nG_91_60 | (nP_91_60 & nG_59_28);
  assign nP_91_28 = nP_91_60 & nP_59_28;
  assign nG_90_27 = nG_90_59 | (nP_90_59 & nG_58_27);
  assign nP_90_27 = nP_90_59 & nP_58_27;
  assign nG_89_26 = nG_89_58 | (nP_89_58 & nG_57_26);
  assign nP_89_26 = nP_89_58 & nP_57_26;
  assign nG_88_25 = nG_88_57 | (nP_88_57 & nG_56_25);
  assign nP_88_25 = nP_88_57 & nP_56_25;
  assign nG_87_24 = nG_87_56 | (nP_87_56 & nG_55_24);
  assign nP_87_24 = nP_87_56 & nP_55_24;
  assign nG_86_23 = nG_86_55 | (nP_86_55 & nG_54_23);
  assign nP_86_23 = nP_86_55 & nP_54_23;
  assign nG_85_22 = nG_85_54 | (nP_85_54 & nG_53_22);
  assign nP_85_22 = nP_85_54 & nP_53_22;
  assign nG_84_21 = nG_84_53 | (nP_84_53 & nG_52_21);
  assign nP_84_21 = nP_84_53 & nP_52_21;
  assign nG_83_20 = nG_83_52 | (nP_83_52 & nG_51_20);
  assign nP_83_20 = nP_83_52 & nP_51_20;
  assign nG_82_19 = nG_82_51 | (nP_82_51 & nG_50_19);
  assign nP_82_19 = nP_82_51 & nP_50_19;
  assign nG_81_18 = nG_81_50 | (nP_81_50 & nG_49_18);
  assign nP_81_18 = nP_81_50 & nP_49_18;
  assign nG_80_17 = nG_80_49 | (nP_80_49 & nG_48_17);
  assign nP_80_17 = nP_80_49 & nP_48_17;
  assign nG_79_16 = nG_79_48 | (nP_79_48 & nG_47_16);
  assign nP_79_16 = nP_79_48 & nP_47_16;
  assign nG_78_15 = nG_78_47 | (nP_78_47 & nG_46_15);
  assign nP_78_15 = nP_78_47 & nP_46_15;
  assign nG_77_14 = nG_77_46 | (nP_77_46 & nG_45_14);
  assign nP_77_14 = nP_77_46 & nP_45_14;
  assign nG_76_13 = nG_76_45 | (nP_76_45 & nG_44_13);
  assign nP_76_13 = nP_76_45 & nP_44_13;
  assign nG_75_12 = nG_75_44 | (nP_75_44 & nG_43_12);
  assign nP_75_12 = nP_75_44 & nP_43_12;
  assign nG_74_11 = nG_74_43 | (nP_74_43 & nG_42_11);
  assign nP_74_11 = nP_74_43 & nP_42_11;
  assign nG_73_10 = nG_73_42 | (nP_73_42 & nG_41_10);
  assign nP_73_10 = nP_73_42 & nP_41_10;
  assign nG_72_9 = nG_72_41 | (nP_72_41 & nG_40_9);
  assign nP_72_9 = nP_72_41 & nP_40_9;
  assign nG_71_8 = nG_71_40 | (nP_71_40 & nG_39_8);
  assign nP_71_8 = nP_71_40 & nP_39_8;
  assign nG_70_7 = nG_70_39 | (nP_70_39 & nG_38_7);
  assign nP_70_7 = nP_70_39 & nP_38_7;
  assign nG_69_6 = nG_69_38 | (nP_69_38 & nG_37_6);
  assign nP_69_6 = nP_69_38 & nP_37_6;
  assign nG_68_5 = nG_68_37 | (nP_68_37 & nG_36_5);
  assign nP_68_5 = nP_68_37 & nP_36_5;
  assign nG_67_4 = nG_67_36 | (nP_67_36 & nG_35_4);
  assign nP_67_4 = nP_67_36 & nP_35_4;
  assign nG_66_3 = nG_66_35 | (nP_66_35 & nG_34_3);
  assign nP_66_3 = nP_66_35 & nP_34_3;
  assign nG_65_2 = nG_65_34 | (nP_65_34 & nG_33_2);
  assign nP_65_2 = nP_65_34 & nP_33_2;
  assign nG_64_1 = nG_64_33 | (nP_64_33 & nG_32_1);
  assign nP_64_1 = nP_64_33 & nP_32_1;
  assign nG_63_0 = nG_63_32 | (nP_63_32 & nG_31_0);
  assign nP_63_0 = nP_63_32 & nP_31_0;
  assign nG_62_0 = nG_62_31 | (nP_62_31 & nG_30_0);
  assign nP_62_0 = nP_62_31 & nP_30_0;
  assign nG_61_0 = nG_61_30 | (nP_61_30 & nG_29_0);
  assign nP_61_0 = nP_61_30 & nP_29_0;
  assign nG_60_0 = nG_60_29 | (nP_60_29 & nG_28_0);
  assign nP_60_0 = nP_60_29 & nP_28_0;
  assign nG_59_0 = nG_59_28 | (nP_59_28 & nG_27_0);
  assign nP_59_0 = nP_59_28 & nP_27_0;
  assign nG_58_0 = nG_58_27 | (nP_58_27 & nG_26_0);
  assign nP_58_0 = nP_58_27 & nP_26_0;
  assign nG_57_0 = nG_57_26 | (nP_57_26 & nG_25_0);
  assign nP_57_0 = nP_57_26 & nP_25_0;
  assign nG_56_0 = nG_56_25 | (nP_56_25 & nG_24_0);
  assign nP_56_0 = nP_56_25 & nP_24_0;
  assign nG_55_0 = nG_55_24 | (nP_55_24 & nG_23_0);
  assign nP_55_0 = nP_55_24 & nP_23_0;
  assign nG_54_0 = nG_54_23 | (nP_54_23 & nG_22_0);
  assign nP_54_0 = nP_54_23 & nP_22_0;
  assign nG_53_0 = nG_53_22 | (nP_53_22 & nG_21_0);
  assign nP_53_0 = nP_53_22 & nP_21_0;
  assign nG_52_0 = nG_52_21 | (nP_52_21 & nG_20_0);
  assign nP_52_0 = nP_52_21 & nP_20_0;
  assign nG_51_0 = nG_51_20 | (nP_51_20 & nG_19_0);
  assign nP_51_0 = nP_51_20 & nP_19_0;
  assign nG_50_0 = nG_50_19 | (nP_50_19 & nG_18_0);
  assign nP_50_0 = nP_50_19 & nP_18_0;
  assign nG_49_0 = nG_49_18 | (nP_49_18 & nG_17_0);
  assign nP_49_0 = nP_49_18 & nP_17_0;
  assign nG_48_0 = nG_48_17 | (nP_48_17 & nG_16_0);
  assign nP_48_0 = nP_48_17 & nP_16_0;
  assign nG_47_0 = nG_47_16 | (nP_47_16 & nG_15_0);
  assign nP_47_0 = nP_47_16 & nP_15_0;
  assign nG_46_0 = nG_46_15 | (nP_46_15 & nG_14_0);
  assign nP_46_0 = nP_46_15 & nP_14_0;
  assign nG_45_0 = nG_45_14 | (nP_45_14 & nG_13_0);
  assign nP_45_0 = nP_45_14 & nP_13_0;
  assign nG_44_0 = nG_44_13 | (nP_44_13 & nG_12_0);
  assign nP_44_0 = nP_44_13 & nP_12_0;
  assign nG_43_0 = nG_43_12 | (nP_43_12 & nG_11_0);
  assign nP_43_0 = nP_43_12 & nP_11_0;
  assign nG_42_0 = nG_42_11 | (nP_42_11 & nG_10_0);
  assign nP_42_0 = nP_42_11 & nP_10_0;
  assign nG_41_0 = nG_41_10 | (nP_41_10 & nG_9_0);
  assign nP_41_0 = nP_41_10 & nP_9_0;
  assign nG_40_0 = nG_40_9 | (nP_40_9 & nG_8_0);
  assign nP_40_0 = nP_40_9 & nP_8_0;
  assign nG_39_0 = nG_39_8 | (nP_39_8 & nG_7_0);
  assign nP_39_0 = nP_39_8 & nP_7_0;
  assign nG_38_0 = nG_38_7 | (nP_38_7 & nG_6_0);
  assign nP_38_0 = nP_38_7 & nP_6_0;
  assign nG_37_0 = nG_37_6 | (nP_37_6 & nG_5_0);
  assign nP_37_0 = nP_37_6 & nP_5_0;
  assign nG_36_0 = nG_36_5 | (nP_36_5 & nG_4_0);
  assign nP_36_0 = nP_36_5 & nP_4_0;
  assign nG_35_0 = nG_35_4 | (nP_35_4 & nG_3_0);
  assign nP_35_0 = nP_35_4 & nP_3_0;
  assign nG_34_0 = nG_34_3 | (nP_34_3 & nG_2_0);
  assign nP_34_0 = nP_34_3 & nP_2_0;
  assign nG_33_0 = nG_33_2 | (nP_33_2 & nG_1_0);
  assign nP_33_0 = nP_33_2 & nP_1_0;
  assign nG_32_0 = nG_32_1 | (nP_32_1 & nG_0_0);
  assign nP_32_0 = nP_32_1 & nP_0_0;

  assign nG_255_128 = nG_255_192 | (nP_255_192 & nG_191_128);
  assign nP_255_128 = nP_255_192 & nP_191_128;
  assign nG_254_127 = nG_254_191 | (nP_254_191 & nG_190_127);
  assign nP_254_127 = nP_254_191 & nP_190_127;
  assign nG_253_126 = nG_253_190 | (nP_253_190 & nG_189_126);
  assign nP_253_126 = nP_253_190 & nP_189_126;
  assign nG_252_125 = nG_252_189 | (nP_252_189 & nG_188_125);
  assign nP_252_125 = nP_252_189 & nP_188_125;
  assign nG_251_124 = nG_251_188 | (nP_251_188 & nG_187_124);
  assign nP_251_124 = nP_251_188 & nP_187_124;
  assign nG_250_123 = nG_250_187 | (nP_250_187 & nG_186_123);
  assign nP_250_123 = nP_250_187 & nP_186_123;
  assign nG_249_122 = nG_249_186 | (nP_249_186 & nG_185_122);
  assign nP_249_122 = nP_249_186 & nP_185_122;
  assign nG_248_121 = nG_248_185 | (nP_248_185 & nG_184_121);
  assign nP_248_121 = nP_248_185 & nP_184_121;
  assign nG_247_120 = nG_247_184 | (nP_247_184 & nG_183_120);
  assign nP_247_120 = nP_247_184 & nP_183_120;
  assign nG_246_119 = nG_246_183 | (nP_246_183 & nG_182_119);
  assign nP_246_119 = nP_246_183 & nP_182_119;
  assign nG_245_118 = nG_245_182 | (nP_245_182 & nG_181_118);
  assign nP_245_118 = nP_245_182 & nP_181_118;
  assign nG_244_117 = nG_244_181 | (nP_244_181 & nG_180_117);
  assign nP_244_117 = nP_244_181 & nP_180_117;
  assign nG_243_116 = nG_243_180 | (nP_243_180 & nG_179_116);
  assign nP_243_116 = nP_243_180 & nP_179_116;
  assign nG_242_115 = nG_242_179 | (nP_242_179 & nG_178_115);
  assign nP_242_115 = nP_242_179 & nP_178_115;
  assign nG_241_114 = nG_241_178 | (nP_241_178 & nG_177_114);
  assign nP_241_114 = nP_241_178 & nP_177_114;
  assign nG_240_113 = nG_240_177 | (nP_240_177 & nG_176_113);
  assign nP_240_113 = nP_240_177 & nP_176_113;
  assign nG_239_112 = nG_239_176 | (nP_239_176 & nG_175_112);
  assign nP_239_112 = nP_239_176 & nP_175_112;
  assign nG_238_111 = nG_238_175 | (nP_238_175 & nG_174_111);
  assign nP_238_111 = nP_238_175 & nP_174_111;
  assign nG_237_110 = nG_237_174 | (nP_237_174 & nG_173_110);
  assign nP_237_110 = nP_237_174 & nP_173_110;
  assign nG_236_109 = nG_236_173 | (nP_236_173 & nG_172_109);
  assign nP_236_109 = nP_236_173 & nP_172_109;
  assign nG_235_108 = nG_235_172 | (nP_235_172 & nG_171_108);
  assign nP_235_108 = nP_235_172 & nP_171_108;
  assign nG_234_107 = nG_234_171 | (nP_234_171 & nG_170_107);
  assign nP_234_107 = nP_234_171 & nP_170_107;
  assign nG_233_106 = nG_233_170 | (nP_233_170 & nG_169_106);
  assign nP_233_106 = nP_233_170 & nP_169_106;
  assign nG_232_105 = nG_232_169 | (nP_232_169 & nG_168_105);
  assign nP_232_105 = nP_232_169 & nP_168_105;
  assign nG_231_104 = nG_231_168 | (nP_231_168 & nG_167_104);
  assign nP_231_104 = nP_231_168 & nP_167_104;
  assign nG_230_103 = nG_230_167 | (nP_230_167 & nG_166_103);
  assign nP_230_103 = nP_230_167 & nP_166_103;
  assign nG_229_102 = nG_229_166 | (nP_229_166 & nG_165_102);
  assign nP_229_102 = nP_229_166 & nP_165_102;
  assign nG_228_101 = nG_228_165 | (nP_228_165 & nG_164_101);
  assign nP_228_101 = nP_228_165 & nP_164_101;
  assign nG_227_100 = nG_227_164 | (nP_227_164 & nG_163_100);
  assign nP_227_100 = nP_227_164 & nP_163_100;
  assign nG_226_99 = nG_226_163 | (nP_226_163 & nG_162_99);
  assign nP_226_99 = nP_226_163 & nP_162_99;
  assign nG_225_98 = nG_225_162 | (nP_225_162 & nG_161_98);
  assign nP_225_98 = nP_225_162 & nP_161_98;
  assign nG_224_97 = nG_224_161 | (nP_224_161 & nG_160_97);
  assign nP_224_97 = nP_224_161 & nP_160_97;
  assign nG_223_96 = nG_223_160 | (nP_223_160 & nG_159_96);
  assign nP_223_96 = nP_223_160 & nP_159_96;
  assign nG_222_95 = nG_222_159 | (nP_222_159 & nG_158_95);
  assign nP_222_95 = nP_222_159 & nP_158_95;
  assign nG_221_94 = nG_221_158 | (nP_221_158 & nG_157_94);
  assign nP_221_94 = nP_221_158 & nP_157_94;
  assign nG_220_93 = nG_220_157 | (nP_220_157 & nG_156_93);
  assign nP_220_93 = nP_220_157 & nP_156_93;
  assign nG_219_92 = nG_219_156 | (nP_219_156 & nG_155_92);
  assign nP_219_92 = nP_219_156 & nP_155_92;
  assign nG_218_91 = nG_218_155 | (nP_218_155 & nG_154_91);
  assign nP_218_91 = nP_218_155 & nP_154_91;
  assign nG_217_90 = nG_217_154 | (nP_217_154 & nG_153_90);
  assign nP_217_90 = nP_217_154 & nP_153_90;
  assign nG_216_89 = nG_216_153 | (nP_216_153 & nG_152_89);
  assign nP_216_89 = nP_216_153 & nP_152_89;
  assign nG_215_88 = nG_215_152 | (nP_215_152 & nG_151_88);
  assign nP_215_88 = nP_215_152 & nP_151_88;
  assign nG_214_87 = nG_214_151 | (nP_214_151 & nG_150_87);
  assign nP_214_87 = nP_214_151 & nP_150_87;
  assign nG_213_86 = nG_213_150 | (nP_213_150 & nG_149_86);
  assign nP_213_86 = nP_213_150 & nP_149_86;
  assign nG_212_85 = nG_212_149 | (nP_212_149 & nG_148_85);
  assign nP_212_85 = nP_212_149 & nP_148_85;
  assign nG_211_84 = nG_211_148 | (nP_211_148 & nG_147_84);
  assign nP_211_84 = nP_211_148 & nP_147_84;
  assign nG_210_83 = nG_210_147 | (nP_210_147 & nG_146_83);
  assign nP_210_83 = nP_210_147 & nP_146_83;
  assign nG_209_82 = nG_209_146 | (nP_209_146 & nG_145_82);
  assign nP_209_82 = nP_209_146 & nP_145_82;
  assign nG_208_81 = nG_208_145 | (nP_208_145 & nG_144_81);
  assign nP_208_81 = nP_208_145 & nP_144_81;
  assign nG_207_80 = nG_207_144 | (nP_207_144 & nG_143_80);
  assign nP_207_80 = nP_207_144 & nP_143_80;
  assign nG_206_79 = nG_206_143 | (nP_206_143 & nG_142_79);
  assign nP_206_79 = nP_206_143 & nP_142_79;
  assign nG_205_78 = nG_205_142 | (nP_205_142 & nG_141_78);
  assign nP_205_78 = nP_205_142 & nP_141_78;
  assign nG_204_77 = nG_204_141 | (nP_204_141 & nG_140_77);
  assign nP_204_77 = nP_204_141 & nP_140_77;
  assign nG_203_76 = nG_203_140 | (nP_203_140 & nG_139_76);
  assign nP_203_76 = nP_203_140 & nP_139_76;
  assign nG_202_75 = nG_202_139 | (nP_202_139 & nG_138_75);
  assign nP_202_75 = nP_202_139 & nP_138_75;
  assign nG_201_74 = nG_201_138 | (nP_201_138 & nG_137_74);
  assign nP_201_74 = nP_201_138 & nP_137_74;
  assign nG_200_73 = nG_200_137 | (nP_200_137 & nG_136_73);
  assign nP_200_73 = nP_200_137 & nP_136_73;
  assign nG_199_72 = nG_199_136 | (nP_199_136 & nG_135_72);
  assign nP_199_72 = nP_199_136 & nP_135_72;
  assign nG_198_71 = nG_198_135 | (nP_198_135 & nG_134_71);
  assign nP_198_71 = nP_198_135 & nP_134_71;
  assign nG_197_70 = nG_197_134 | (nP_197_134 & nG_133_70);
  assign nP_197_70 = nP_197_134 & nP_133_70;
  assign nG_196_69 = nG_196_133 | (nP_196_133 & nG_132_69);
  assign nP_196_69 = nP_196_133 & nP_132_69;
  assign nG_195_68 = nG_195_132 | (nP_195_132 & nG_131_68);
  assign nP_195_68 = nP_195_132 & nP_131_68;
  assign nG_194_67 = nG_194_131 | (nP_194_131 & nG_130_67);
  assign nP_194_67 = nP_194_131 & nP_130_67;
  assign nG_193_66 = nG_193_130 | (nP_193_130 & nG_129_66);
  assign nP_193_66 = nP_193_130 & nP_129_66;
  assign nG_192_65 = nG_192_129 | (nP_192_129 & nG_128_65);
  assign nP_192_65 = nP_192_129 & nP_128_65;
  assign nG_191_64 = nG_191_128 | (nP_191_128 & nG_127_64);
  assign nP_191_64 = nP_191_128 & nP_127_64;
  assign nG_190_63 = nG_190_127 | (nP_190_127 & nG_126_63);
  assign nP_190_63 = nP_190_127 & nP_126_63;
  assign nG_189_62 = nG_189_126 | (nP_189_126 & nG_125_62);
  assign nP_189_62 = nP_189_126 & nP_125_62;
  assign nG_188_61 = nG_188_125 | (nP_188_125 & nG_124_61);
  assign nP_188_61 = nP_188_125 & nP_124_61;
  assign nG_187_60 = nG_187_124 | (nP_187_124 & nG_123_60);
  assign nP_187_60 = nP_187_124 & nP_123_60;
  assign nG_186_59 = nG_186_123 | (nP_186_123 & nG_122_59);
  assign nP_186_59 = nP_186_123 & nP_122_59;
  assign nG_185_58 = nG_185_122 | (nP_185_122 & nG_121_58);
  assign nP_185_58 = nP_185_122 & nP_121_58;
  assign nG_184_57 = nG_184_121 | (nP_184_121 & nG_120_57);
  assign nP_184_57 = nP_184_121 & nP_120_57;
  assign nG_183_56 = nG_183_120 | (nP_183_120 & nG_119_56);
  assign nP_183_56 = nP_183_120 & nP_119_56;
  assign nG_182_55 = nG_182_119 | (nP_182_119 & nG_118_55);
  assign nP_182_55 = nP_182_119 & nP_118_55;
  assign nG_181_54 = nG_181_118 | (nP_181_118 & nG_117_54);
  assign nP_181_54 = nP_181_118 & nP_117_54;
  assign nG_180_53 = nG_180_117 | (nP_180_117 & nG_116_53);
  assign nP_180_53 = nP_180_117 & nP_116_53;
  assign nG_179_52 = nG_179_116 | (nP_179_116 & nG_115_52);
  assign nP_179_52 = nP_179_116 & nP_115_52;
  assign nG_178_51 = nG_178_115 | (nP_178_115 & nG_114_51);
  assign nP_178_51 = nP_178_115 & nP_114_51;
  assign nG_177_50 = nG_177_114 | (nP_177_114 & nG_113_50);
  assign nP_177_50 = nP_177_114 & nP_113_50;
  assign nG_176_49 = nG_176_113 | (nP_176_113 & nG_112_49);
  assign nP_176_49 = nP_176_113 & nP_112_49;
  assign nG_175_48 = nG_175_112 | (nP_175_112 & nG_111_48);
  assign nP_175_48 = nP_175_112 & nP_111_48;
  assign nG_174_47 = nG_174_111 | (nP_174_111 & nG_110_47);
  assign nP_174_47 = nP_174_111 & nP_110_47;
  assign nG_173_46 = nG_173_110 | (nP_173_110 & nG_109_46);
  assign nP_173_46 = nP_173_110 & nP_109_46;
  assign nG_172_45 = nG_172_109 | (nP_172_109 & nG_108_45);
  assign nP_172_45 = nP_172_109 & nP_108_45;
  assign nG_171_44 = nG_171_108 | (nP_171_108 & nG_107_44);
  assign nP_171_44 = nP_171_108 & nP_107_44;
  assign nG_170_43 = nG_170_107 | (nP_170_107 & nG_106_43);
  assign nP_170_43 = nP_170_107 & nP_106_43;
  assign nG_169_42 = nG_169_106 | (nP_169_106 & nG_105_42);
  assign nP_169_42 = nP_169_106 & nP_105_42;
  assign nG_168_41 = nG_168_105 | (nP_168_105 & nG_104_41);
  assign nP_168_41 = nP_168_105 & nP_104_41;
  assign nG_167_40 = nG_167_104 | (nP_167_104 & nG_103_40);
  assign nP_167_40 = nP_167_104 & nP_103_40;
  assign nG_166_39 = nG_166_103 | (nP_166_103 & nG_102_39);
  assign nP_166_39 = nP_166_103 & nP_102_39;
  assign nG_165_38 = nG_165_102 | (nP_165_102 & nG_101_38);
  assign nP_165_38 = nP_165_102 & nP_101_38;
  assign nG_164_37 = nG_164_101 | (nP_164_101 & nG_100_37);
  assign nP_164_37 = nP_164_101 & nP_100_37;
  assign nG_163_36 = nG_163_100 | (nP_163_100 & nG_99_36);
  assign nP_163_36 = nP_163_100 & nP_99_36;
  assign nG_162_35 = nG_162_99 | (nP_162_99 & nG_98_35);
  assign nP_162_35 = nP_162_99 & nP_98_35;
  assign nG_161_34 = nG_161_98 | (nP_161_98 & nG_97_34);
  assign nP_161_34 = nP_161_98 & nP_97_34;
  assign nG_160_33 = nG_160_97 | (nP_160_97 & nG_96_33);
  assign nP_160_33 = nP_160_97 & nP_96_33;
  assign nG_159_32 = nG_159_96 | (nP_159_96 & nG_95_32);
  assign nP_159_32 = nP_159_96 & nP_95_32;
  assign nG_158_31 = nG_158_95 | (nP_158_95 & nG_94_31);
  assign nP_158_31 = nP_158_95 & nP_94_31;
  assign nG_157_30 = nG_157_94 | (nP_157_94 & nG_93_30);
  assign nP_157_30 = nP_157_94 & nP_93_30;
  assign nG_156_29 = nG_156_93 | (nP_156_93 & nG_92_29);
  assign nP_156_29 = nP_156_93 & nP_92_29;
  assign nG_155_28 = nG_155_92 | (nP_155_92 & nG_91_28);
  assign nP_155_28 = nP_155_92 & nP_91_28;
  assign nG_154_27 = nG_154_91 | (nP_154_91 & nG_90_27);
  assign nP_154_27 = nP_154_91 & nP_90_27;
  assign nG_153_26 = nG_153_90 | (nP_153_90 & nG_89_26);
  assign nP_153_26 = nP_153_90 & nP_89_26;
  assign nG_152_25 = nG_152_89 | (nP_152_89 & nG_88_25);
  assign nP_152_25 = nP_152_89 & nP_88_25;
  assign nG_151_24 = nG_151_88 | (nP_151_88 & nG_87_24);
  assign nP_151_24 = nP_151_88 & nP_87_24;
  assign nG_150_23 = nG_150_87 | (nP_150_87 & nG_86_23);
  assign nP_150_23 = nP_150_87 & nP_86_23;
  assign nG_149_22 = nG_149_86 | (nP_149_86 & nG_85_22);
  assign nP_149_22 = nP_149_86 & nP_85_22;
  assign nG_148_21 = nG_148_85 | (nP_148_85 & nG_84_21);
  assign nP_148_21 = nP_148_85 & nP_84_21;
  assign nG_147_20 = nG_147_84 | (nP_147_84 & nG_83_20);
  assign nP_147_20 = nP_147_84 & nP_83_20;
  assign nG_146_19 = nG_146_83 | (nP_146_83 & nG_82_19);
  assign nP_146_19 = nP_146_83 & nP_82_19;
  assign nG_145_18 = nG_145_82 | (nP_145_82 & nG_81_18);
  assign nP_145_18 = nP_145_82 & nP_81_18;
  assign nG_144_17 = nG_144_81 | (nP_144_81 & nG_80_17);
  assign nP_144_17 = nP_144_81 & nP_80_17;
  assign nG_143_16 = nG_143_80 | (nP_143_80 & nG_79_16);
  assign nP_143_16 = nP_143_80 & nP_79_16;
  assign nG_142_15 = nG_142_79 | (nP_142_79 & nG_78_15);
  assign nP_142_15 = nP_142_79 & nP_78_15;
  assign nG_141_14 = nG_141_78 | (nP_141_78 & nG_77_14);
  assign nP_141_14 = nP_141_78 & nP_77_14;
  assign nG_140_13 = nG_140_77 | (nP_140_77 & nG_76_13);
  assign nP_140_13 = nP_140_77 & nP_76_13;
  assign nG_139_12 = nG_139_76 | (nP_139_76 & nG_75_12);
  assign nP_139_12 = nP_139_76 & nP_75_12;
  assign nG_138_11 = nG_138_75 | (nP_138_75 & nG_74_11);
  assign nP_138_11 = nP_138_75 & nP_74_11;
  assign nG_137_10 = nG_137_74 | (nP_137_74 & nG_73_10);
  assign nP_137_10 = nP_137_74 & nP_73_10;
  assign nG_136_9 = nG_136_73 | (nP_136_73 & nG_72_9);
  assign nP_136_9 = nP_136_73 & nP_72_9;
  assign nG_135_8 = nG_135_72 | (nP_135_72 & nG_71_8);
  assign nP_135_8 = nP_135_72 & nP_71_8;
  assign nG_134_7 = nG_134_71 | (nP_134_71 & nG_70_7);
  assign nP_134_7 = nP_134_71 & nP_70_7;
  assign nG_133_6 = nG_133_70 | (nP_133_70 & nG_69_6);
  assign nP_133_6 = nP_133_70 & nP_69_6;
  assign nG_132_5 = nG_132_69 | (nP_132_69 & nG_68_5);
  assign nP_132_5 = nP_132_69 & nP_68_5;
  assign nG_131_4 = nG_131_68 | (nP_131_68 & nG_67_4);
  assign nP_131_4 = nP_131_68 & nP_67_4;
  assign nG_130_3 = nG_130_67 | (nP_130_67 & nG_66_3);
  assign nP_130_3 = nP_130_67 & nP_66_3;
  assign nG_129_2 = nG_129_66 | (nP_129_66 & nG_65_2);
  assign nP_129_2 = nP_129_66 & nP_65_2;
  assign nG_128_1 = nG_128_65 | (nP_128_65 & nG_64_1);
  assign nP_128_1 = nP_128_65 & nP_64_1;
  assign nG_127_0 = nG_127_64 | (nP_127_64 & nG_63_0);
  assign nP_127_0 = nP_127_64 & nP_63_0;
  assign nG_126_0 = nG_126_63 | (nP_126_63 & nG_62_0);
  assign nP_126_0 = nP_126_63 & nP_62_0;
  assign nG_125_0 = nG_125_62 | (nP_125_62 & nG_61_0);
  assign nP_125_0 = nP_125_62 & nP_61_0;
  assign nG_124_0 = nG_124_61 | (nP_124_61 & nG_60_0);
  assign nP_124_0 = nP_124_61 & nP_60_0;
  assign nG_123_0 = nG_123_60 | (nP_123_60 & nG_59_0);
  assign nP_123_0 = nP_123_60 & nP_59_0;
  assign nG_122_0 = nG_122_59 | (nP_122_59 & nG_58_0);
  assign nP_122_0 = nP_122_59 & nP_58_0;
  assign nG_121_0 = nG_121_58 | (nP_121_58 & nG_57_0);
  assign nP_121_0 = nP_121_58 & nP_57_0;
  assign nG_120_0 = nG_120_57 | (nP_120_57 & nG_56_0);
  assign nP_120_0 = nP_120_57 & nP_56_0;
  assign nG_119_0 = nG_119_56 | (nP_119_56 & nG_55_0);
  assign nP_119_0 = nP_119_56 & nP_55_0;
  assign nG_118_0 = nG_118_55 | (nP_118_55 & nG_54_0);
  assign nP_118_0 = nP_118_55 & nP_54_0;
  assign nG_117_0 = nG_117_54 | (nP_117_54 & nG_53_0);
  assign nP_117_0 = nP_117_54 & nP_53_0;
  assign nG_116_0 = nG_116_53 | (nP_116_53 & nG_52_0);
  assign nP_116_0 = nP_116_53 & nP_52_0;
  assign nG_115_0 = nG_115_52 | (nP_115_52 & nG_51_0);
  assign nP_115_0 = nP_115_52 & nP_51_0;
  assign nG_114_0 = nG_114_51 | (nP_114_51 & nG_50_0);
  assign nP_114_0 = nP_114_51 & nP_50_0;
  assign nG_113_0 = nG_113_50 | (nP_113_50 & nG_49_0);
  assign nP_113_0 = nP_113_50 & nP_49_0;
  assign nG_112_0 = nG_112_49 | (nP_112_49 & nG_48_0);
  assign nP_112_0 = nP_112_49 & nP_48_0;
  assign nG_111_0 = nG_111_48 | (nP_111_48 & nG_47_0);
  assign nP_111_0 = nP_111_48 & nP_47_0;
  assign nG_110_0 = nG_110_47 | (nP_110_47 & nG_46_0);
  assign nP_110_0 = nP_110_47 & nP_46_0;
  assign nG_109_0 = nG_109_46 | (nP_109_46 & nG_45_0);
  assign nP_109_0 = nP_109_46 & nP_45_0;
  assign nG_108_0 = nG_108_45 | (nP_108_45 & nG_44_0);
  assign nP_108_0 = nP_108_45 & nP_44_0;
  assign nG_107_0 = nG_107_44 | (nP_107_44 & nG_43_0);
  assign nP_107_0 = nP_107_44 & nP_43_0;
  assign nG_106_0 = nG_106_43 | (nP_106_43 & nG_42_0);
  assign nP_106_0 = nP_106_43 & nP_42_0;
  assign nG_105_0 = nG_105_42 | (nP_105_42 & nG_41_0);
  assign nP_105_0 = nP_105_42 & nP_41_0;
  assign nG_104_0 = nG_104_41 | (nP_104_41 & nG_40_0);
  assign nP_104_0 = nP_104_41 & nP_40_0;
  assign nG_103_0 = nG_103_40 | (nP_103_40 & nG_39_0);
  assign nP_103_0 = nP_103_40 & nP_39_0;
  assign nG_102_0 = nG_102_39 | (nP_102_39 & nG_38_0);
  assign nP_102_0 = nP_102_39 & nP_38_0;
  assign nG_101_0 = nG_101_38 | (nP_101_38 & nG_37_0);
  assign nP_101_0 = nP_101_38 & nP_37_0;
  assign nG_100_0 = nG_100_37 | (nP_100_37 & nG_36_0);
  assign nP_100_0 = nP_100_37 & nP_36_0;
  assign nG_99_0 = nG_99_36 | (nP_99_36 & nG_35_0);
  assign nP_99_0 = nP_99_36 & nP_35_0;
  assign nG_98_0 = nG_98_35 | (nP_98_35 & nG_34_0);
  assign nP_98_0 = nP_98_35 & nP_34_0;
  assign nG_97_0 = nG_97_34 | (nP_97_34 & nG_33_0);
  assign nP_97_0 = nP_97_34 & nP_33_0;
  assign nG_96_0 = nG_96_33 | (nP_96_33 & nG_32_0);
  assign nP_96_0 = nP_96_33 & nP_32_0;
  assign nG_95_0 = nG_95_32 | (nP_95_32 & nG_31_0);
  assign nP_95_0 = nP_95_32 & nP_31_0;
  assign nG_94_0 = nG_94_31 | (nP_94_31 & nG_30_0);
  assign nP_94_0 = nP_94_31 & nP_30_0;
  assign nG_93_0 = nG_93_30 | (nP_93_30 & nG_29_0);
  assign nP_93_0 = nP_93_30 & nP_29_0;
  assign nG_92_0 = nG_92_29 | (nP_92_29 & nG_28_0);
  assign nP_92_0 = nP_92_29 & nP_28_0;
  assign nG_91_0 = nG_91_28 | (nP_91_28 & nG_27_0);
  assign nP_91_0 = nP_91_28 & nP_27_0;
  assign nG_90_0 = nG_90_27 | (nP_90_27 & nG_26_0);
  assign nP_90_0 = nP_90_27 & nP_26_0;
  assign nG_89_0 = nG_89_26 | (nP_89_26 & nG_25_0);
  assign nP_89_0 = nP_89_26 & nP_25_0;
  assign nG_88_0 = nG_88_25 | (nP_88_25 & nG_24_0);
  assign nP_88_0 = nP_88_25 & nP_24_0;
  assign nG_87_0 = nG_87_24 | (nP_87_24 & nG_23_0);
  assign nP_87_0 = nP_87_24 & nP_23_0;
  assign nG_86_0 = nG_86_23 | (nP_86_23 & nG_22_0);
  assign nP_86_0 = nP_86_23 & nP_22_0;
  assign nG_85_0 = nG_85_22 | (nP_85_22 & nG_21_0);
  assign nP_85_0 = nP_85_22 & nP_21_0;
  assign nG_84_0 = nG_84_21 | (nP_84_21 & nG_20_0);
  assign nP_84_0 = nP_84_21 & nP_20_0;
  assign nG_83_0 = nG_83_20 | (nP_83_20 & nG_19_0);
  assign nP_83_0 = nP_83_20 & nP_19_0;
  assign nG_82_0 = nG_82_19 | (nP_82_19 & nG_18_0);
  assign nP_82_0 = nP_82_19 & nP_18_0;
  assign nG_81_0 = nG_81_18 | (nP_81_18 & nG_17_0);
  assign nP_81_0 = nP_81_18 & nP_17_0;
  assign nG_80_0 = nG_80_17 | (nP_80_17 & nG_16_0);
  assign nP_80_0 = nP_80_17 & nP_16_0;
  assign nG_79_0 = nG_79_16 | (nP_79_16 & nG_15_0);
  assign nP_79_0 = nP_79_16 & nP_15_0;
  assign nG_78_0 = nG_78_15 | (nP_78_15 & nG_14_0);
  assign nP_78_0 = nP_78_15 & nP_14_0;
  assign nG_77_0 = nG_77_14 | (nP_77_14 & nG_13_0);
  assign nP_77_0 = nP_77_14 & nP_13_0;
  assign nG_76_0 = nG_76_13 | (nP_76_13 & nG_12_0);
  assign nP_76_0 = nP_76_13 & nP_12_0;
  assign nG_75_0 = nG_75_12 | (nP_75_12 & nG_11_0);
  assign nP_75_0 = nP_75_12 & nP_11_0;
  assign nG_74_0 = nG_74_11 | (nP_74_11 & nG_10_0);
  assign nP_74_0 = nP_74_11 & nP_10_0;
  assign nG_73_0 = nG_73_10 | (nP_73_10 & nG_9_0);
  assign nP_73_0 = nP_73_10 & nP_9_0;
  assign nG_72_0 = nG_72_9 | (nP_72_9 & nG_8_0);
  assign nP_72_0 = nP_72_9 & nP_8_0;
  assign nG_71_0 = nG_71_8 | (nP_71_8 & nG_7_0);
  assign nP_71_0 = nP_71_8 & nP_7_0;
  assign nG_70_0 = nG_70_7 | (nP_70_7 & nG_6_0);
  assign nP_70_0 = nP_70_7 & nP_6_0;
  assign nG_69_0 = nG_69_6 | (nP_69_6 & nG_5_0);
  assign nP_69_0 = nP_69_6 & nP_5_0;
  assign nG_68_0 = nG_68_5 | (nP_68_5 & nG_4_0);
  assign nP_68_0 = nP_68_5 & nP_4_0;
  assign nG_67_0 = nG_67_4 | (nP_67_4 & nG_3_0);
  assign nP_67_0 = nP_67_4 & nP_3_0;
  assign nG_66_0 = nG_66_3 | (nP_66_3 & nG_2_0);
  assign nP_66_0 = nP_66_3 & nP_2_0;
  assign nG_65_0 = nG_65_2 | (nP_65_2 & nG_1_0);
  assign nP_65_0 = nP_65_2 & nP_1_0;
  assign nG_64_0 = nG_64_1 | (nP_64_1 & nG_0_0);
  assign nP_64_0 = nP_64_1 & nP_0_0;

  assign nG_255_0 = nG_255_128 | (nP_255_128 & nG_127_0);
  assign nP_255_0 = nP_255_128 & nP_127_0;
  assign nG_254_0 = nG_254_127 | (nP_254_127 & nG_126_0);
  assign nP_254_0 = nP_254_127 & nP_126_0;
  assign nG_253_0 = nG_253_126 | (nP_253_126 & nG_125_0);
  assign nP_253_0 = nP_253_126 & nP_125_0;
  assign nG_252_0 = nG_252_125 | (nP_252_125 & nG_124_0);
  assign nP_252_0 = nP_252_125 & nP_124_0;
  assign nG_251_0 = nG_251_124 | (nP_251_124 & nG_123_0);
  assign nP_251_0 = nP_251_124 & nP_123_0;
  assign nG_250_0 = nG_250_123 | (nP_250_123 & nG_122_0);
  assign nP_250_0 = nP_250_123 & nP_122_0;
  assign nG_249_0 = nG_249_122 | (nP_249_122 & nG_121_0);
  assign nP_249_0 = nP_249_122 & nP_121_0;
  assign nG_248_0 = nG_248_121 | (nP_248_121 & nG_120_0);
  assign nP_248_0 = nP_248_121 & nP_120_0;
  assign nG_247_0 = nG_247_120 | (nP_247_120 & nG_119_0);
  assign nP_247_0 = nP_247_120 & nP_119_0;
  assign nG_246_0 = nG_246_119 | (nP_246_119 & nG_118_0);
  assign nP_246_0 = nP_246_119 & nP_118_0;
  assign nG_245_0 = nG_245_118 | (nP_245_118 & nG_117_0);
  assign nP_245_0 = nP_245_118 & nP_117_0;
  assign nG_244_0 = nG_244_117 | (nP_244_117 & nG_116_0);
  assign nP_244_0 = nP_244_117 & nP_116_0;
  assign nG_243_0 = nG_243_116 | (nP_243_116 & nG_115_0);
  assign nP_243_0 = nP_243_116 & nP_115_0;
  assign nG_242_0 = nG_242_115 | (nP_242_115 & nG_114_0);
  assign nP_242_0 = nP_242_115 & nP_114_0;
  assign nG_241_0 = nG_241_114 | (nP_241_114 & nG_113_0);
  assign nP_241_0 = nP_241_114 & nP_113_0;
  assign nG_240_0 = nG_240_113 | (nP_240_113 & nG_112_0);
  assign nP_240_0 = nP_240_113 & nP_112_0;
  assign nG_239_0 = nG_239_112 | (nP_239_112 & nG_111_0);
  assign nP_239_0 = nP_239_112 & nP_111_0;
  assign nG_238_0 = nG_238_111 | (nP_238_111 & nG_110_0);
  assign nP_238_0 = nP_238_111 & nP_110_0;
  assign nG_237_0 = nG_237_110 | (nP_237_110 & nG_109_0);
  assign nP_237_0 = nP_237_110 & nP_109_0;
  assign nG_236_0 = nG_236_109 | (nP_236_109 & nG_108_0);
  assign nP_236_0 = nP_236_109 & nP_108_0;
  assign nG_235_0 = nG_235_108 | (nP_235_108 & nG_107_0);
  assign nP_235_0 = nP_235_108 & nP_107_0;
  assign nG_234_0 = nG_234_107 | (nP_234_107 & nG_106_0);
  assign nP_234_0 = nP_234_107 & nP_106_0;
  assign nG_233_0 = nG_233_106 | (nP_233_106 & nG_105_0);
  assign nP_233_0 = nP_233_106 & nP_105_0;
  assign nG_232_0 = nG_232_105 | (nP_232_105 & nG_104_0);
  assign nP_232_0 = nP_232_105 & nP_104_0;
  assign nG_231_0 = nG_231_104 | (nP_231_104 & nG_103_0);
  assign nP_231_0 = nP_231_104 & nP_103_0;
  assign nG_230_0 = nG_230_103 | (nP_230_103 & nG_102_0);
  assign nP_230_0 = nP_230_103 & nP_102_0;
  assign nG_229_0 = nG_229_102 | (nP_229_102 & nG_101_0);
  assign nP_229_0 = nP_229_102 & nP_101_0;
  assign nG_228_0 = nG_228_101 | (nP_228_101 & nG_100_0);
  assign nP_228_0 = nP_228_101 & nP_100_0;
  assign nG_227_0 = nG_227_100 | (nP_227_100 & nG_99_0);
  assign nP_227_0 = nP_227_100 & nP_99_0;
  assign nG_226_0 = nG_226_99 | (nP_226_99 & nG_98_0);
  assign nP_226_0 = nP_226_99 & nP_98_0;
  assign nG_225_0 = nG_225_98 | (nP_225_98 & nG_97_0);
  assign nP_225_0 = nP_225_98 & nP_97_0;
  assign nG_224_0 = nG_224_97 | (nP_224_97 & nG_96_0);
  assign nP_224_0 = nP_224_97 & nP_96_0;
  assign nG_223_0 = nG_223_96 | (nP_223_96 & nG_95_0);
  assign nP_223_0 = nP_223_96 & nP_95_0;
  assign nG_222_0 = nG_222_95 | (nP_222_95 & nG_94_0);
  assign nP_222_0 = nP_222_95 & nP_94_0;
  assign nG_221_0 = nG_221_94 | (nP_221_94 & nG_93_0);
  assign nP_221_0 = nP_221_94 & nP_93_0;
  assign nG_220_0 = nG_220_93 | (nP_220_93 & nG_92_0);
  assign nP_220_0 = nP_220_93 & nP_92_0;
  assign nG_219_0 = nG_219_92 | (nP_219_92 & nG_91_0);
  assign nP_219_0 = nP_219_92 & nP_91_0;
  assign nG_218_0 = nG_218_91 | (nP_218_91 & nG_90_0);
  assign nP_218_0 = nP_218_91 & nP_90_0;
  assign nG_217_0 = nG_217_90 | (nP_217_90 & nG_89_0);
  assign nP_217_0 = nP_217_90 & nP_89_0;
  assign nG_216_0 = nG_216_89 | (nP_216_89 & nG_88_0);
  assign nP_216_0 = nP_216_89 & nP_88_0;
  assign nG_215_0 = nG_215_88 | (nP_215_88 & nG_87_0);
  assign nP_215_0 = nP_215_88 & nP_87_0;
  assign nG_214_0 = nG_214_87 | (nP_214_87 & nG_86_0);
  assign nP_214_0 = nP_214_87 & nP_86_0;
  assign nG_213_0 = nG_213_86 | (nP_213_86 & nG_85_0);
  assign nP_213_0 = nP_213_86 & nP_85_0;
  assign nG_212_0 = nG_212_85 | (nP_212_85 & nG_84_0);
  assign nP_212_0 = nP_212_85 & nP_84_0;
  assign nG_211_0 = nG_211_84 | (nP_211_84 & nG_83_0);
  assign nP_211_0 = nP_211_84 & nP_83_0;
  assign nG_210_0 = nG_210_83 | (nP_210_83 & nG_82_0);
  assign nP_210_0 = nP_210_83 & nP_82_0;
  assign nG_209_0 = nG_209_82 | (nP_209_82 & nG_81_0);
  assign nP_209_0 = nP_209_82 & nP_81_0;
  assign nG_208_0 = nG_208_81 | (nP_208_81 & nG_80_0);
  assign nP_208_0 = nP_208_81 & nP_80_0;
  assign nG_207_0 = nG_207_80 | (nP_207_80 & nG_79_0);
  assign nP_207_0 = nP_207_80 & nP_79_0;
  assign nG_206_0 = nG_206_79 | (nP_206_79 & nG_78_0);
  assign nP_206_0 = nP_206_79 & nP_78_0;
  assign nG_205_0 = nG_205_78 | (nP_205_78 & nG_77_0);
  assign nP_205_0 = nP_205_78 & nP_77_0;
  assign nG_204_0 = nG_204_77 | (nP_204_77 & nG_76_0);
  assign nP_204_0 = nP_204_77 & nP_76_0;
  assign nG_203_0 = nG_203_76 | (nP_203_76 & nG_75_0);
  assign nP_203_0 = nP_203_76 & nP_75_0;
  assign nG_202_0 = nG_202_75 | (nP_202_75 & nG_74_0);
  assign nP_202_0 = nP_202_75 & nP_74_0;
  assign nG_201_0 = nG_201_74 | (nP_201_74 & nG_73_0);
  assign nP_201_0 = nP_201_74 & nP_73_0;
  assign nG_200_0 = nG_200_73 | (nP_200_73 & nG_72_0);
  assign nP_200_0 = nP_200_73 & nP_72_0;
  assign nG_199_0 = nG_199_72 | (nP_199_72 & nG_71_0);
  assign nP_199_0 = nP_199_72 & nP_71_0;
  assign nG_198_0 = nG_198_71 | (nP_198_71 & nG_70_0);
  assign nP_198_0 = nP_198_71 & nP_70_0;
  assign nG_197_0 = nG_197_70 | (nP_197_70 & nG_69_0);
  assign nP_197_0 = nP_197_70 & nP_69_0;
  assign nG_196_0 = nG_196_69 | (nP_196_69 & nG_68_0);
  assign nP_196_0 = nP_196_69 & nP_68_0;
  assign nG_195_0 = nG_195_68 | (nP_195_68 & nG_67_0);
  assign nP_195_0 = nP_195_68 & nP_67_0;
  assign nG_194_0 = nG_194_67 | (nP_194_67 & nG_66_0);
  assign nP_194_0 = nP_194_67 & nP_66_0;
  assign nG_193_0 = nG_193_66 | (nP_193_66 & nG_65_0);
  assign nP_193_0 = nP_193_66 & nP_65_0;
  assign nG_192_0 = nG_192_65 | (nP_192_65 & nG_64_0);
  assign nP_192_0 = nP_192_65 & nP_64_0;
  assign nG_191_0 = nG_191_64 | (nP_191_64 & nG_63_0);
  assign nP_191_0 = nP_191_64 & nP_63_0;
  assign nG_190_0 = nG_190_63 | (nP_190_63 & nG_62_0);
  assign nP_190_0 = nP_190_63 & nP_62_0;
  assign nG_189_0 = nG_189_62 | (nP_189_62 & nG_61_0);
  assign nP_189_0 = nP_189_62 & nP_61_0;
  assign nG_188_0 = nG_188_61 | (nP_188_61 & nG_60_0);
  assign nP_188_0 = nP_188_61 & nP_60_0;
  assign nG_187_0 = nG_187_60 | (nP_187_60 & nG_59_0);
  assign nP_187_0 = nP_187_60 & nP_59_0;
  assign nG_186_0 = nG_186_59 | (nP_186_59 & nG_58_0);
  assign nP_186_0 = nP_186_59 & nP_58_0;
  assign nG_185_0 = nG_185_58 | (nP_185_58 & nG_57_0);
  assign nP_185_0 = nP_185_58 & nP_57_0;
  assign nG_184_0 = nG_184_57 | (nP_184_57 & nG_56_0);
  assign nP_184_0 = nP_184_57 & nP_56_0;
  assign nG_183_0 = nG_183_56 | (nP_183_56 & nG_55_0);
  assign nP_183_0 = nP_183_56 & nP_55_0;
  assign nG_182_0 = nG_182_55 | (nP_182_55 & nG_54_0);
  assign nP_182_0 = nP_182_55 & nP_54_0;
  assign nG_181_0 = nG_181_54 | (nP_181_54 & nG_53_0);
  assign nP_181_0 = nP_181_54 & nP_53_0;
  assign nG_180_0 = nG_180_53 | (nP_180_53 & nG_52_0);
  assign nP_180_0 = nP_180_53 & nP_52_0;
  assign nG_179_0 = nG_179_52 | (nP_179_52 & nG_51_0);
  assign nP_179_0 = nP_179_52 & nP_51_0;
  assign nG_178_0 = nG_178_51 | (nP_178_51 & nG_50_0);
  assign nP_178_0 = nP_178_51 & nP_50_0;
  assign nG_177_0 = nG_177_50 | (nP_177_50 & nG_49_0);
  assign nP_177_0 = nP_177_50 & nP_49_0;
  assign nG_176_0 = nG_176_49 | (nP_176_49 & nG_48_0);
  assign nP_176_0 = nP_176_49 & nP_48_0;
  assign nG_175_0 = nG_175_48 | (nP_175_48 & nG_47_0);
  assign nP_175_0 = nP_175_48 & nP_47_0;
  assign nG_174_0 = nG_174_47 | (nP_174_47 & nG_46_0);
  assign nP_174_0 = nP_174_47 & nP_46_0;
  assign nG_173_0 = nG_173_46 | (nP_173_46 & nG_45_0);
  assign nP_173_0 = nP_173_46 & nP_45_0;
  assign nG_172_0 = nG_172_45 | (nP_172_45 & nG_44_0);
  assign nP_172_0 = nP_172_45 & nP_44_0;
  assign nG_171_0 = nG_171_44 | (nP_171_44 & nG_43_0);
  assign nP_171_0 = nP_171_44 & nP_43_0;
  assign nG_170_0 = nG_170_43 | (nP_170_43 & nG_42_0);
  assign nP_170_0 = nP_170_43 & nP_42_0;
  assign nG_169_0 = nG_169_42 | (nP_169_42 & nG_41_0);
  assign nP_169_0 = nP_169_42 & nP_41_0;
  assign nG_168_0 = nG_168_41 | (nP_168_41 & nG_40_0);
  assign nP_168_0 = nP_168_41 & nP_40_0;
  assign nG_167_0 = nG_167_40 | (nP_167_40 & nG_39_0);
  assign nP_167_0 = nP_167_40 & nP_39_0;
  assign nG_166_0 = nG_166_39 | (nP_166_39 & nG_38_0);
  assign nP_166_0 = nP_166_39 & nP_38_0;
  assign nG_165_0 = nG_165_38 | (nP_165_38 & nG_37_0);
  assign nP_165_0 = nP_165_38 & nP_37_0;
  assign nG_164_0 = nG_164_37 | (nP_164_37 & nG_36_0);
  assign nP_164_0 = nP_164_37 & nP_36_0;
  assign nG_163_0 = nG_163_36 | (nP_163_36 & nG_35_0);
  assign nP_163_0 = nP_163_36 & nP_35_0;
  assign nG_162_0 = nG_162_35 | (nP_162_35 & nG_34_0);
  assign nP_162_0 = nP_162_35 & nP_34_0;
  assign nG_161_0 = nG_161_34 | (nP_161_34 & nG_33_0);
  assign nP_161_0 = nP_161_34 & nP_33_0;
  assign nG_160_0 = nG_160_33 | (nP_160_33 & nG_32_0);
  assign nP_160_0 = nP_160_33 & nP_32_0;
  assign nG_159_0 = nG_159_32 | (nP_159_32 & nG_31_0);
  assign nP_159_0 = nP_159_32 & nP_31_0;
  assign nG_158_0 = nG_158_31 | (nP_158_31 & nG_30_0);
  assign nP_158_0 = nP_158_31 & nP_30_0;
  assign nG_157_0 = nG_157_30 | (nP_157_30 & nG_29_0);
  assign nP_157_0 = nP_157_30 & nP_29_0;
  assign nG_156_0 = nG_156_29 | (nP_156_29 & nG_28_0);
  assign nP_156_0 = nP_156_29 & nP_28_0;
  assign nG_155_0 = nG_155_28 | (nP_155_28 & nG_27_0);
  assign nP_155_0 = nP_155_28 & nP_27_0;
  assign nG_154_0 = nG_154_27 | (nP_154_27 & nG_26_0);
  assign nP_154_0 = nP_154_27 & nP_26_0;
  assign nG_153_0 = nG_153_26 | (nP_153_26 & nG_25_0);
  assign nP_153_0 = nP_153_26 & nP_25_0;
  assign nG_152_0 = nG_152_25 | (nP_152_25 & nG_24_0);
  assign nP_152_0 = nP_152_25 & nP_24_0;
  assign nG_151_0 = nG_151_24 | (nP_151_24 & nG_23_0);
  assign nP_151_0 = nP_151_24 & nP_23_0;
  assign nG_150_0 = nG_150_23 | (nP_150_23 & nG_22_0);
  assign nP_150_0 = nP_150_23 & nP_22_0;
  assign nG_149_0 = nG_149_22 | (nP_149_22 & nG_21_0);
  assign nP_149_0 = nP_149_22 & nP_21_0;
  assign nG_148_0 = nG_148_21 | (nP_148_21 & nG_20_0);
  assign nP_148_0 = nP_148_21 & nP_20_0;
  assign nG_147_0 = nG_147_20 | (nP_147_20 & nG_19_0);
  assign nP_147_0 = nP_147_20 & nP_19_0;
  assign nG_146_0 = nG_146_19 | (nP_146_19 & nG_18_0);
  assign nP_146_0 = nP_146_19 & nP_18_0;
  assign nG_145_0 = nG_145_18 | (nP_145_18 & nG_17_0);
  assign nP_145_0 = nP_145_18 & nP_17_0;
  assign nG_144_0 = nG_144_17 | (nP_144_17 & nG_16_0);
  assign nP_144_0 = nP_144_17 & nP_16_0;
  assign nG_143_0 = nG_143_16 | (nP_143_16 & nG_15_0);
  assign nP_143_0 = nP_143_16 & nP_15_0;
  assign nG_142_0 = nG_142_15 | (nP_142_15 & nG_14_0);
  assign nP_142_0 = nP_142_15 & nP_14_0;
  assign nG_141_0 = nG_141_14 | (nP_141_14 & nG_13_0);
  assign nP_141_0 = nP_141_14 & nP_13_0;
  assign nG_140_0 = nG_140_13 | (nP_140_13 & nG_12_0);
  assign nP_140_0 = nP_140_13 & nP_12_0;
  assign nG_139_0 = nG_139_12 | (nP_139_12 & nG_11_0);
  assign nP_139_0 = nP_139_12 & nP_11_0;
  assign nG_138_0 = nG_138_11 | (nP_138_11 & nG_10_0);
  assign nP_138_0 = nP_138_11 & nP_10_0;
  assign nG_137_0 = nG_137_10 | (nP_137_10 & nG_9_0);
  assign nP_137_0 = nP_137_10 & nP_9_0;
  assign nG_136_0 = nG_136_9 | (nP_136_9 & nG_8_0);
  assign nP_136_0 = nP_136_9 & nP_8_0;
  assign nG_135_0 = nG_135_8 | (nP_135_8 & nG_7_0);
  assign nP_135_0 = nP_135_8 & nP_7_0;
  assign nG_134_0 = nG_134_7 | (nP_134_7 & nG_6_0);
  assign nP_134_0 = nP_134_7 & nP_6_0;
  assign nG_133_0 = nG_133_6 | (nP_133_6 & nG_5_0);
  assign nP_133_0 = nP_133_6 & nP_5_0;
  assign nG_132_0 = nG_132_5 | (nP_132_5 & nG_4_0);
  assign nP_132_0 = nP_132_5 & nP_4_0;
  assign nG_131_0 = nG_131_4 | (nP_131_4 & nG_3_0);
  assign nP_131_0 = nP_131_4 & nP_3_0;
  assign nG_130_0 = nG_130_3 | (nP_130_3 & nG_2_0);
  assign nP_130_0 = nP_130_3 & nP_2_0;
  assign nG_129_0 = nG_129_2 | (nP_129_2 & nG_1_0);
  assign nP_129_0 = nP_129_2 & nP_1_0;
  assign nG_128_0 = nG_128_1 | (nP_128_1 & nG_0_0);
  assign nP_128_0 = nP_128_1 & nP_0_0;

  assign nC_0 = in_CI;
  assign nC_1 = nG_0_0 | (nP_0_0 & in_CI);
  assign nC_2 = nG_1_0 | (nP_1_0 & in_CI);
  assign nC_3 = nG_2_0 | (nP_2_0 & in_CI);
  assign nC_4 = nG_3_0 | (nP_3_0 & in_CI);
  assign nC_5 = nG_4_0 | (nP_4_0 & in_CI);
  assign nC_6 = nG_5_0 | (nP_5_0 & in_CI);
  assign nC_7 = nG_6_0 | (nP_6_0 & in_CI);
  assign nC_8 = nG_7_0 | (nP_7_0 & in_CI);
  assign nC_9 = nG_8_0 | (nP_8_0 & in_CI);
  assign nC_10 = nG_9_0 | (nP_9_0 & in_CI);
  assign nC_11 = nG_10_0 | (nP_10_0 & in_CI);
  assign nC_12 = nG_11_0 | (nP_11_0 & in_CI);
  assign nC_13 = nG_12_0 | (nP_12_0 & in_CI);
  assign nC_14 = nG_13_0 | (nP_13_0 & in_CI);
  assign nC_15 = nG_14_0 | (nP_14_0 & in_CI);
  assign nC_16 = nG_15_0 | (nP_15_0 & in_CI);
  assign nC_17 = nG_16_0 | (nP_16_0 & in_CI);
  assign nC_18 = nG_17_0 | (nP_17_0 & in_CI);
  assign nC_19 = nG_18_0 | (nP_18_0 & in_CI);
  assign nC_20 = nG_19_0 | (nP_19_0 & in_CI);
  assign nC_21 = nG_20_0 | (nP_20_0 & in_CI);
  assign nC_22 = nG_21_0 | (nP_21_0 & in_CI);
  assign nC_23 = nG_22_0 | (nP_22_0 & in_CI);
  assign nC_24 = nG_23_0 | (nP_23_0 & in_CI);
  assign nC_25 = nG_24_0 | (nP_24_0 & in_CI);
  assign nC_26 = nG_25_0 | (nP_25_0 & in_CI);
  assign nC_27 = nG_26_0 | (nP_26_0 & in_CI);
  assign nC_28 = nG_27_0 | (nP_27_0 & in_CI);
  assign nC_29 = nG_28_0 | (nP_28_0 & in_CI);
  assign nC_30 = nG_29_0 | (nP_29_0 & in_CI);
  assign nC_31 = nG_30_0 | (nP_30_0 & in_CI);
  assign nC_32 = nG_31_0 | (nP_31_0 & in_CI);
  assign nC_33 = nG_32_0 | (nP_32_0 & in_CI);
  assign nC_34 = nG_33_0 | (nP_33_0 & in_CI);
  assign nC_35 = nG_34_0 | (nP_34_0 & in_CI);
  assign nC_36 = nG_35_0 | (nP_35_0 & in_CI);
  assign nC_37 = nG_36_0 | (nP_36_0 & in_CI);
  assign nC_38 = nG_37_0 | (nP_37_0 & in_CI);
  assign nC_39 = nG_38_0 | (nP_38_0 & in_CI);
  assign nC_40 = nG_39_0 | (nP_39_0 & in_CI);
  assign nC_41 = nG_40_0 | (nP_40_0 & in_CI);
  assign nC_42 = nG_41_0 | (nP_41_0 & in_CI);
  assign nC_43 = nG_42_0 | (nP_42_0 & in_CI);
  assign nC_44 = nG_43_0 | (nP_43_0 & in_CI);
  assign nC_45 = nG_44_0 | (nP_44_0 & in_CI);
  assign nC_46 = nG_45_0 | (nP_45_0 & in_CI);
  assign nC_47 = nG_46_0 | (nP_46_0 & in_CI);
  assign nC_48 = nG_47_0 | (nP_47_0 & in_CI);
  assign nC_49 = nG_48_0 | (nP_48_0 & in_CI);
  assign nC_50 = nG_49_0 | (nP_49_0 & in_CI);
  assign nC_51 = nG_50_0 | (nP_50_0 & in_CI);
  assign nC_52 = nG_51_0 | (nP_51_0 & in_CI);
  assign nC_53 = nG_52_0 | (nP_52_0 & in_CI);
  assign nC_54 = nG_53_0 | (nP_53_0 & in_CI);
  assign nC_55 = nG_54_0 | (nP_54_0 & in_CI);
  assign nC_56 = nG_55_0 | (nP_55_0 & in_CI);
  assign nC_57 = nG_56_0 | (nP_56_0 & in_CI);
  assign nC_58 = nG_57_0 | (nP_57_0 & in_CI);
  assign nC_59 = nG_58_0 | (nP_58_0 & in_CI);
  assign nC_60 = nG_59_0 | (nP_59_0 & in_CI);
  assign nC_61 = nG_60_0 | (nP_60_0 & in_CI);
  assign nC_62 = nG_61_0 | (nP_61_0 & in_CI);
  assign nC_63 = nG_62_0 | (nP_62_0 & in_CI);
  assign nC_64 = nG_63_0 | (nP_63_0 & in_CI);
  assign nC_65 = nG_64_0 | (nP_64_0 & in_CI);
  assign nC_66 = nG_65_0 | (nP_65_0 & in_CI);
  assign nC_67 = nG_66_0 | (nP_66_0 & in_CI);
  assign nC_68 = nG_67_0 | (nP_67_0 & in_CI);
  assign nC_69 = nG_68_0 | (nP_68_0 & in_CI);
  assign nC_70 = nG_69_0 | (nP_69_0 & in_CI);
  assign nC_71 = nG_70_0 | (nP_70_0 & in_CI);
  assign nC_72 = nG_71_0 | (nP_71_0 & in_CI);
  assign nC_73 = nG_72_0 | (nP_72_0 & in_CI);
  assign nC_74 = nG_73_0 | (nP_73_0 & in_CI);
  assign nC_75 = nG_74_0 | (nP_74_0 & in_CI);
  assign nC_76 = nG_75_0 | (nP_75_0 & in_CI);
  assign nC_77 = nG_76_0 | (nP_76_0 & in_CI);
  assign nC_78 = nG_77_0 | (nP_77_0 & in_CI);
  assign nC_79 = nG_78_0 | (nP_78_0 & in_CI);
  assign nC_80 = nG_79_0 | (nP_79_0 & in_CI);
  assign nC_81 = nG_80_0 | (nP_80_0 & in_CI);
  assign nC_82 = nG_81_0 | (nP_81_0 & in_CI);
  assign nC_83 = nG_82_0 | (nP_82_0 & in_CI);
  assign nC_84 = nG_83_0 | (nP_83_0 & in_CI);
  assign nC_85 = nG_84_0 | (nP_84_0 & in_CI);
  assign nC_86 = nG_85_0 | (nP_85_0 & in_CI);
  assign nC_87 = nG_86_0 | (nP_86_0 & in_CI);
  assign nC_88 = nG_87_0 | (nP_87_0 & in_CI);
  assign nC_89 = nG_88_0 | (nP_88_0 & in_CI);
  assign nC_90 = nG_89_0 | (nP_89_0 & in_CI);
  assign nC_91 = nG_90_0 | (nP_90_0 & in_CI);
  assign nC_92 = nG_91_0 | (nP_91_0 & in_CI);
  assign nC_93 = nG_92_0 | (nP_92_0 & in_CI);
  assign nC_94 = nG_93_0 | (nP_93_0 & in_CI);
  assign nC_95 = nG_94_0 | (nP_94_0 & in_CI);
  assign nC_96 = nG_95_0 | (nP_95_0 & in_CI);
  assign nC_97 = nG_96_0 | (nP_96_0 & in_CI);
  assign nC_98 = nG_97_0 | (nP_97_0 & in_CI);
  assign nC_99 = nG_98_0 | (nP_98_0 & in_CI);
  assign nC_100 = nG_99_0 | (nP_99_0 & in_CI);
  assign nC_101 = nG_100_0 | (nP_100_0 & in_CI);
  assign nC_102 = nG_101_0 | (nP_101_0 & in_CI);
  assign nC_103 = nG_102_0 | (nP_102_0 & in_CI);
  assign nC_104 = nG_103_0 | (nP_103_0 & in_CI);
  assign nC_105 = nG_104_0 | (nP_104_0 & in_CI);
  assign nC_106 = nG_105_0 | (nP_105_0 & in_CI);
  assign nC_107 = nG_106_0 | (nP_106_0 & in_CI);
  assign nC_108 = nG_107_0 | (nP_107_0 & in_CI);
  assign nC_109 = nG_108_0 | (nP_108_0 & in_CI);
  assign nC_110 = nG_109_0 | (nP_109_0 & in_CI);
  assign nC_111 = nG_110_0 | (nP_110_0 & in_CI);
  assign nC_112 = nG_111_0 | (nP_111_0 & in_CI);
  assign nC_113 = nG_112_0 | (nP_112_0 & in_CI);
  assign nC_114 = nG_113_0 | (nP_113_0 & in_CI);
  assign nC_115 = nG_114_0 | (nP_114_0 & in_CI);
  assign nC_116 = nG_115_0 | (nP_115_0 & in_CI);
  assign nC_117 = nG_116_0 | (nP_116_0 & in_CI);
  assign nC_118 = nG_117_0 | (nP_117_0 & in_CI);
  assign nC_119 = nG_118_0 | (nP_118_0 & in_CI);
  assign nC_120 = nG_119_0 | (nP_119_0 & in_CI);
  assign nC_121 = nG_120_0 | (nP_120_0 & in_CI);
  assign nC_122 = nG_121_0 | (nP_121_0 & in_CI);
  assign nC_123 = nG_122_0 | (nP_122_0 & in_CI);
  assign nC_124 = nG_123_0 | (nP_123_0 & in_CI);
  assign nC_125 = nG_124_0 | (nP_124_0 & in_CI);
  assign nC_126 = nG_125_0 | (nP_125_0 & in_CI);
  assign nC_127 = nG_126_0 | (nP_126_0 & in_CI);
  assign nC_128 = nG_127_0 | (nP_127_0 & in_CI);
  assign nC_129 = nG_128_0 | (nP_128_0 & in_CI);
  assign nC_130 = nG_129_0 | (nP_129_0 & in_CI);
  assign nC_131 = nG_130_0 | (nP_130_0 & in_CI);
  assign nC_132 = nG_131_0 | (nP_131_0 & in_CI);
  assign nC_133 = nG_132_0 | (nP_132_0 & in_CI);
  assign nC_134 = nG_133_0 | (nP_133_0 & in_CI);
  assign nC_135 = nG_134_0 | (nP_134_0 & in_CI);
  assign nC_136 = nG_135_0 | (nP_135_0 & in_CI);
  assign nC_137 = nG_136_0 | (nP_136_0 & in_CI);
  assign nC_138 = nG_137_0 | (nP_137_0 & in_CI);
  assign nC_139 = nG_138_0 | (nP_138_0 & in_CI);
  assign nC_140 = nG_139_0 | (nP_139_0 & in_CI);
  assign nC_141 = nG_140_0 | (nP_140_0 & in_CI);
  assign nC_142 = nG_141_0 | (nP_141_0 & in_CI);
  assign nC_143 = nG_142_0 | (nP_142_0 & in_CI);
  assign nC_144 = nG_143_0 | (nP_143_0 & in_CI);
  assign nC_145 = nG_144_0 | (nP_144_0 & in_CI);
  assign nC_146 = nG_145_0 | (nP_145_0 & in_CI);
  assign nC_147 = nG_146_0 | (nP_146_0 & in_CI);
  assign nC_148 = nG_147_0 | (nP_147_0 & in_CI);
  assign nC_149 = nG_148_0 | (nP_148_0 & in_CI);
  assign nC_150 = nG_149_0 | (nP_149_0 & in_CI);
  assign nC_151 = nG_150_0 | (nP_150_0 & in_CI);
  assign nC_152 = nG_151_0 | (nP_151_0 & in_CI);
  assign nC_153 = nG_152_0 | (nP_152_0 & in_CI);
  assign nC_154 = nG_153_0 | (nP_153_0 & in_CI);
  assign nC_155 = nG_154_0 | (nP_154_0 & in_CI);
  assign nC_156 = nG_155_0 | (nP_155_0 & in_CI);
  assign nC_157 = nG_156_0 | (nP_156_0 & in_CI);
  assign nC_158 = nG_157_0 | (nP_157_0 & in_CI);
  assign nC_159 = nG_158_0 | (nP_158_0 & in_CI);
  assign nC_160 = nG_159_0 | (nP_159_0 & in_CI);
  assign nC_161 = nG_160_0 | (nP_160_0 & in_CI);
  assign nC_162 = nG_161_0 | (nP_161_0 & in_CI);
  assign nC_163 = nG_162_0 | (nP_162_0 & in_CI);
  assign nC_164 = nG_163_0 | (nP_163_0 & in_CI);
  assign nC_165 = nG_164_0 | (nP_164_0 & in_CI);
  assign nC_166 = nG_165_0 | (nP_165_0 & in_CI);
  assign nC_167 = nG_166_0 | (nP_166_0 & in_CI);
  assign nC_168 = nG_167_0 | (nP_167_0 & in_CI);
  assign nC_169 = nG_168_0 | (nP_168_0 & in_CI);
  assign nC_170 = nG_169_0 | (nP_169_0 & in_CI);
  assign nC_171 = nG_170_0 | (nP_170_0 & in_CI);
  assign nC_172 = nG_171_0 | (nP_171_0 & in_CI);
  assign nC_173 = nG_172_0 | (nP_172_0 & in_CI);
  assign nC_174 = nG_173_0 | (nP_173_0 & in_CI);
  assign nC_175 = nG_174_0 | (nP_174_0 & in_CI);
  assign nC_176 = nG_175_0 | (nP_175_0 & in_CI);
  assign nC_177 = nG_176_0 | (nP_176_0 & in_CI);
  assign nC_178 = nG_177_0 | (nP_177_0 & in_CI);
  assign nC_179 = nG_178_0 | (nP_178_0 & in_CI);
  assign nC_180 = nG_179_0 | (nP_179_0 & in_CI);
  assign nC_181 = nG_180_0 | (nP_180_0 & in_CI);
  assign nC_182 = nG_181_0 | (nP_181_0 & in_CI);
  assign nC_183 = nG_182_0 | (nP_182_0 & in_CI);
  assign nC_184 = nG_183_0 | (nP_183_0 & in_CI);
  assign nC_185 = nG_184_0 | (nP_184_0 & in_CI);
  assign nC_186 = nG_185_0 | (nP_185_0 & in_CI);
  assign nC_187 = nG_186_0 | (nP_186_0 & in_CI);
  assign nC_188 = nG_187_0 | (nP_187_0 & in_CI);
  assign nC_189 = nG_188_0 | (nP_188_0 & in_CI);
  assign nC_190 = nG_189_0 | (nP_189_0 & in_CI);
  assign nC_191 = nG_190_0 | (nP_190_0 & in_CI);
  assign nC_192 = nG_191_0 | (nP_191_0 & in_CI);
  assign nC_193 = nG_192_0 | (nP_192_0 & in_CI);
  assign nC_194 = nG_193_0 | (nP_193_0 & in_CI);
  assign nC_195 = nG_194_0 | (nP_194_0 & in_CI);
  assign nC_196 = nG_195_0 | (nP_195_0 & in_CI);
  assign nC_197 = nG_196_0 | (nP_196_0 & in_CI);
  assign nC_198 = nG_197_0 | (nP_197_0 & in_CI);
  assign nC_199 = nG_198_0 | (nP_198_0 & in_CI);
  assign nC_200 = nG_199_0 | (nP_199_0 & in_CI);
  assign nC_201 = nG_200_0 | (nP_200_0 & in_CI);
  assign nC_202 = nG_201_0 | (nP_201_0 & in_CI);
  assign nC_203 = nG_202_0 | (nP_202_0 & in_CI);
  assign nC_204 = nG_203_0 | (nP_203_0 & in_CI);
  assign nC_205 = nG_204_0 | (nP_204_0 & in_CI);
  assign nC_206 = nG_205_0 | (nP_205_0 & in_CI);
  assign nC_207 = nG_206_0 | (nP_206_0 & in_CI);
  assign nC_208 = nG_207_0 | (nP_207_0 & in_CI);
  assign nC_209 = nG_208_0 | (nP_208_0 & in_CI);
  assign nC_210 = nG_209_0 | (nP_209_0 & in_CI);
  assign nC_211 = nG_210_0 | (nP_210_0 & in_CI);
  assign nC_212 = nG_211_0 | (nP_211_0 & in_CI);
  assign nC_213 = nG_212_0 | (nP_212_0 & in_CI);
  assign nC_214 = nG_213_0 | (nP_213_0 & in_CI);
  assign nC_215 = nG_214_0 | (nP_214_0 & in_CI);
  assign nC_216 = nG_215_0 | (nP_215_0 & in_CI);
  assign nC_217 = nG_216_0 | (nP_216_0 & in_CI);
  assign nC_218 = nG_217_0 | (nP_217_0 & in_CI);
  assign nC_219 = nG_218_0 | (nP_218_0 & in_CI);
  assign nC_220 = nG_219_0 | (nP_219_0 & in_CI);
  assign nC_221 = nG_220_0 | (nP_220_0 & in_CI);
  assign nC_222 = nG_221_0 | (nP_221_0 & in_CI);
  assign nC_223 = nG_222_0 | (nP_222_0 & in_CI);
  assign nC_224 = nG_223_0 | (nP_223_0 & in_CI);
  assign nC_225 = nG_224_0 | (nP_224_0 & in_CI);
  assign nC_226 = nG_225_0 | (nP_225_0 & in_CI);
  assign nC_227 = nG_226_0 | (nP_226_0 & in_CI);
  assign nC_228 = nG_227_0 | (nP_227_0 & in_CI);
  assign nC_229 = nG_228_0 | (nP_228_0 & in_CI);
  assign nC_230 = nG_229_0 | (nP_229_0 & in_CI);
  assign nC_231 = nG_230_0 | (nP_230_0 & in_CI);
  assign nC_232 = nG_231_0 | (nP_231_0 & in_CI);
  assign nC_233 = nG_232_0 | (nP_232_0 & in_CI);
  assign nC_234 = nG_233_0 | (nP_233_0 & in_CI);
  assign nC_235 = nG_234_0 | (nP_234_0 & in_CI);
  assign nC_236 = nG_235_0 | (nP_235_0 & in_CI);
  assign nC_237 = nG_236_0 | (nP_236_0 & in_CI);
  assign nC_238 = nG_237_0 | (nP_237_0 & in_CI);
  assign nC_239 = nG_238_0 | (nP_238_0 & in_CI);
  assign nC_240 = nG_239_0 | (nP_239_0 & in_CI);
  assign nC_241 = nG_240_0 | (nP_240_0 & in_CI);
  assign nC_242 = nG_241_0 | (nP_241_0 & in_CI);
  assign nC_243 = nG_242_0 | (nP_242_0 & in_CI);
  assign nC_244 = nG_243_0 | (nP_243_0 & in_CI);
  assign nC_245 = nG_244_0 | (nP_244_0 & in_CI);
  assign nC_246 = nG_245_0 | (nP_245_0 & in_CI);
  assign nC_247 = nG_246_0 | (nP_246_0 & in_CI);
  assign nC_248 = nG_247_0 | (nP_247_0 & in_CI);
  assign nC_249 = nG_248_0 | (nP_248_0 & in_CI);
  assign nC_250 = nG_249_0 | (nP_249_0 & in_CI);
  assign nC_251 = nG_250_0 | (nP_250_0 & in_CI);
  assign nC_252 = nG_251_0 | (nP_251_0 & in_CI);
  assign nC_253 = nG_252_0 | (nP_252_0 & in_CI);
  assign nC_254 = nG_253_0 | (nP_253_0 & in_CI);
  assign nC_255 = nG_254_0 | (nP_254_0 & in_CI);

  assign out_S[0] = nP_0_0 ^ nC_0;
  assign out_S[1] = nP_1_1 ^ nC_1;
  assign out_S[2] = nP_2_2 ^ nC_2;
  assign out_S[3] = nP_3_3 ^ nC_3;
  assign out_S[4] = nP_4_4 ^ nC_4;
  assign out_S[5] = nP_5_5 ^ nC_5;
  assign out_S[6] = nP_6_6 ^ nC_6;
  assign out_S[7] = nP_7_7 ^ nC_7;
  assign out_S[8] = nP_8_8 ^ nC_8;
  assign out_S[9] = nP_9_9 ^ nC_9;
  assign out_S[10] = nP_10_10 ^ nC_10;
  assign out_S[11] = nP_11_11 ^ nC_11;
  assign out_S[12] = nP_12_12 ^ nC_12;
  assign out_S[13] = nP_13_13 ^ nC_13;
  assign out_S[14] = nP_14_14 ^ nC_14;
  assign out_S[15] = nP_15_15 ^ nC_15;
  assign out_S[16] = nP_16_16 ^ nC_16;
  assign out_S[17] = nP_17_17 ^ nC_17;
  assign out_S[18] = nP_18_18 ^ nC_18;
  assign out_S[19] = nP_19_19 ^ nC_19;
  assign out_S[20] = nP_20_20 ^ nC_20;
  assign out_S[21] = nP_21_21 ^ nC_21;
  assign out_S[22] = nP_22_22 ^ nC_22;
  assign out_S[23] = nP_23_23 ^ nC_23;
  assign out_S[24] = nP_24_24 ^ nC_24;
  assign out_S[25] = nP_25_25 ^ nC_25;
  assign out_S[26] = nP_26_26 ^ nC_26;
  assign out_S[27] = nP_27_27 ^ nC_27;
  assign out_S[28] = nP_28_28 ^ nC_28;
  assign out_S[29] = nP_29_29 ^ nC_29;
  assign out_S[30] = nP_30_30 ^ nC_30;
  assign out_S[31] = nP_31_31 ^ nC_31;
  assign out_S[32] = nP_32_32 ^ nC_32;
  assign out_S[33] = nP_33_33 ^ nC_33;
  assign out_S[34] = nP_34_34 ^ nC_34;
  assign out_S[35] = nP_35_35 ^ nC_35;
  assign out_S[36] = nP_36_36 ^ nC_36;
  assign out_S[37] = nP_37_37 ^ nC_37;
  assign out_S[38] = nP_38_38 ^ nC_38;
  assign out_S[39] = nP_39_39 ^ nC_39;
  assign out_S[40] = nP_40_40 ^ nC_40;
  assign out_S[41] = nP_41_41 ^ nC_41;
  assign out_S[42] = nP_42_42 ^ nC_42;
  assign out_S[43] = nP_43_43 ^ nC_43;
  assign out_S[44] = nP_44_44 ^ nC_44;
  assign out_S[45] = nP_45_45 ^ nC_45;
  assign out_S[46] = nP_46_46 ^ nC_46;
  assign out_S[47] = nP_47_47 ^ nC_47;
  assign out_S[48] = nP_48_48 ^ nC_48;
  assign out_S[49] = nP_49_49 ^ nC_49;
  assign out_S[50] = nP_50_50 ^ nC_50;
  assign out_S[51] = nP_51_51 ^ nC_51;
  assign out_S[52] = nP_52_52 ^ nC_52;
  assign out_S[53] = nP_53_53 ^ nC_53;
  assign out_S[54] = nP_54_54 ^ nC_54;
  assign out_S[55] = nP_55_55 ^ nC_55;
  assign out_S[56] = nP_56_56 ^ nC_56;
  assign out_S[57] = nP_57_57 ^ nC_57;
  assign out_S[58] = nP_58_58 ^ nC_58;
  assign out_S[59] = nP_59_59 ^ nC_59;
  assign out_S[60] = nP_60_60 ^ nC_60;
  assign out_S[61] = nP_61_61 ^ nC_61;
  assign out_S[62] = nP_62_62 ^ nC_62;
  assign out_S[63] = nP_63_63 ^ nC_63;
  assign out_S[64] = nP_64_64 ^ nC_64;
  assign out_S[65] = nP_65_65 ^ nC_65;
  assign out_S[66] = nP_66_66 ^ nC_66;
  assign out_S[67] = nP_67_67 ^ nC_67;
  assign out_S[68] = nP_68_68 ^ nC_68;
  assign out_S[69] = nP_69_69 ^ nC_69;
  assign out_S[70] = nP_70_70 ^ nC_70;
  assign out_S[71] = nP_71_71 ^ nC_71;
  assign out_S[72] = nP_72_72 ^ nC_72;
  assign out_S[73] = nP_73_73 ^ nC_73;
  assign out_S[74] = nP_74_74 ^ nC_74;
  assign out_S[75] = nP_75_75 ^ nC_75;
  assign out_S[76] = nP_76_76 ^ nC_76;
  assign out_S[77] = nP_77_77 ^ nC_77;
  assign out_S[78] = nP_78_78 ^ nC_78;
  assign out_S[79] = nP_79_79 ^ nC_79;
  assign out_S[80] = nP_80_80 ^ nC_80;
  assign out_S[81] = nP_81_81 ^ nC_81;
  assign out_S[82] = nP_82_82 ^ nC_82;
  assign out_S[83] = nP_83_83 ^ nC_83;
  assign out_S[84] = nP_84_84 ^ nC_84;
  assign out_S[85] = nP_85_85 ^ nC_85;
  assign out_S[86] = nP_86_86 ^ nC_86;
  assign out_S[87] = nP_87_87 ^ nC_87;
  assign out_S[88] = nP_88_88 ^ nC_88;
  assign out_S[89] = nP_89_89 ^ nC_89;
  assign out_S[90] = nP_90_90 ^ nC_90;
  assign out_S[91] = nP_91_91 ^ nC_91;
  assign out_S[92] = nP_92_92 ^ nC_92;
  assign out_S[93] = nP_93_93 ^ nC_93;
  assign out_S[94] = nP_94_94 ^ nC_94;
  assign out_S[95] = nP_95_95 ^ nC_95;
  assign out_S[96] = nP_96_96 ^ nC_96;
  assign out_S[97] = nP_97_97 ^ nC_97;
  assign out_S[98] = nP_98_98 ^ nC_98;
  assign out_S[99] = nP_99_99 ^ nC_99;
  assign out_S[100] = nP_100_100 ^ nC_100;
  assign out_S[101] = nP_101_101 ^ nC_101;
  assign out_S[102] = nP_102_102 ^ nC_102;
  assign out_S[103] = nP_103_103 ^ nC_103;
  assign out_S[104] = nP_104_104 ^ nC_104;
  assign out_S[105] = nP_105_105 ^ nC_105;
  assign out_S[106] = nP_106_106 ^ nC_106;
  assign out_S[107] = nP_107_107 ^ nC_107;
  assign out_S[108] = nP_108_108 ^ nC_108;
  assign out_S[109] = nP_109_109 ^ nC_109;
  assign out_S[110] = nP_110_110 ^ nC_110;
  assign out_S[111] = nP_111_111 ^ nC_111;
  assign out_S[112] = nP_112_112 ^ nC_112;
  assign out_S[113] = nP_113_113 ^ nC_113;
  assign out_S[114] = nP_114_114 ^ nC_114;
  assign out_S[115] = nP_115_115 ^ nC_115;
  assign out_S[116] = nP_116_116 ^ nC_116;
  assign out_S[117] = nP_117_117 ^ nC_117;
  assign out_S[118] = nP_118_118 ^ nC_118;
  assign out_S[119] = nP_119_119 ^ nC_119;
  assign out_S[120] = nP_120_120 ^ nC_120;
  assign out_S[121] = nP_121_121 ^ nC_121;
  assign out_S[122] = nP_122_122 ^ nC_122;
  assign out_S[123] = nP_123_123 ^ nC_123;
  assign out_S[124] = nP_124_124 ^ nC_124;
  assign out_S[125] = nP_125_125 ^ nC_125;
  assign out_S[126] = nP_126_126 ^ nC_126;
  assign out_S[127] = nP_127_127 ^ nC_127;
  assign out_S[128] = nP_128_128 ^ nC_128;
  assign out_S[129] = nP_129_129 ^ nC_129;
  assign out_S[130] = nP_130_130 ^ nC_130;
  assign out_S[131] = nP_131_131 ^ nC_131;
  assign out_S[132] = nP_132_132 ^ nC_132;
  assign out_S[133] = nP_133_133 ^ nC_133;
  assign out_S[134] = nP_134_134 ^ nC_134;
  assign out_S[135] = nP_135_135 ^ nC_135;
  assign out_S[136] = nP_136_136 ^ nC_136;
  assign out_S[137] = nP_137_137 ^ nC_137;
  assign out_S[138] = nP_138_138 ^ nC_138;
  assign out_S[139] = nP_139_139 ^ nC_139;
  assign out_S[140] = nP_140_140 ^ nC_140;
  assign out_S[141] = nP_141_141 ^ nC_141;
  assign out_S[142] = nP_142_142 ^ nC_142;
  assign out_S[143] = nP_143_143 ^ nC_143;
  assign out_S[144] = nP_144_144 ^ nC_144;
  assign out_S[145] = nP_145_145 ^ nC_145;
  assign out_S[146] = nP_146_146 ^ nC_146;
  assign out_S[147] = nP_147_147 ^ nC_147;
  assign out_S[148] = nP_148_148 ^ nC_148;
  assign out_S[149] = nP_149_149 ^ nC_149;
  assign out_S[150] = nP_150_150 ^ nC_150;
  assign out_S[151] = nP_151_151 ^ nC_151;
  assign out_S[152] = nP_152_152 ^ nC_152;
  assign out_S[153] = nP_153_153 ^ nC_153;
  assign out_S[154] = nP_154_154 ^ nC_154;
  assign out_S[155] = nP_155_155 ^ nC_155;
  assign out_S[156] = nP_156_156 ^ nC_156;
  assign out_S[157] = nP_157_157 ^ nC_157;
  assign out_S[158] = nP_158_158 ^ nC_158;
  assign out_S[159] = nP_159_159 ^ nC_159;
  assign out_S[160] = nP_160_160 ^ nC_160;
  assign out_S[161] = nP_161_161 ^ nC_161;
  assign out_S[162] = nP_162_162 ^ nC_162;
  assign out_S[163] = nP_163_163 ^ nC_163;
  assign out_S[164] = nP_164_164 ^ nC_164;
  assign out_S[165] = nP_165_165 ^ nC_165;
  assign out_S[166] = nP_166_166 ^ nC_166;
  assign out_S[167] = nP_167_167 ^ nC_167;
  assign out_S[168] = nP_168_168 ^ nC_168;
  assign out_S[169] = nP_169_169 ^ nC_169;
  assign out_S[170] = nP_170_170 ^ nC_170;
  assign out_S[171] = nP_171_171 ^ nC_171;
  assign out_S[172] = nP_172_172 ^ nC_172;
  assign out_S[173] = nP_173_173 ^ nC_173;
  assign out_S[174] = nP_174_174 ^ nC_174;
  assign out_S[175] = nP_175_175 ^ nC_175;
  assign out_S[176] = nP_176_176 ^ nC_176;
  assign out_S[177] = nP_177_177 ^ nC_177;
  assign out_S[178] = nP_178_178 ^ nC_178;
  assign out_S[179] = nP_179_179 ^ nC_179;
  assign out_S[180] = nP_180_180 ^ nC_180;
  assign out_S[181] = nP_181_181 ^ nC_181;
  assign out_S[182] = nP_182_182 ^ nC_182;
  assign out_S[183] = nP_183_183 ^ nC_183;
  assign out_S[184] = nP_184_184 ^ nC_184;
  assign out_S[185] = nP_185_185 ^ nC_185;
  assign out_S[186] = nP_186_186 ^ nC_186;
  assign out_S[187] = nP_187_187 ^ nC_187;
  assign out_S[188] = nP_188_188 ^ nC_188;
  assign out_S[189] = nP_189_189 ^ nC_189;
  assign out_S[190] = nP_190_190 ^ nC_190;
  assign out_S[191] = nP_191_191 ^ nC_191;
  assign out_S[192] = nP_192_192 ^ nC_192;
  assign out_S[193] = nP_193_193 ^ nC_193;
  assign out_S[194] = nP_194_194 ^ nC_194;
  assign out_S[195] = nP_195_195 ^ nC_195;
  assign out_S[196] = nP_196_196 ^ nC_196;
  assign out_S[197] = nP_197_197 ^ nC_197;
  assign out_S[198] = nP_198_198 ^ nC_198;
  assign out_S[199] = nP_199_199 ^ nC_199;
  assign out_S[200] = nP_200_200 ^ nC_200;
  assign out_S[201] = nP_201_201 ^ nC_201;
  assign out_S[202] = nP_202_202 ^ nC_202;
  assign out_S[203] = nP_203_203 ^ nC_203;
  assign out_S[204] = nP_204_204 ^ nC_204;
  assign out_S[205] = nP_205_205 ^ nC_205;
  assign out_S[206] = nP_206_206 ^ nC_206;
  assign out_S[207] = nP_207_207 ^ nC_207;
  assign out_S[208] = nP_208_208 ^ nC_208;
  assign out_S[209] = nP_209_209 ^ nC_209;
  assign out_S[210] = nP_210_210 ^ nC_210;
  assign out_S[211] = nP_211_211 ^ nC_211;
  assign out_S[212] = nP_212_212 ^ nC_212;
  assign out_S[213] = nP_213_213 ^ nC_213;
  assign out_S[214] = nP_214_214 ^ nC_214;
  assign out_S[215] = nP_215_215 ^ nC_215;
  assign out_S[216] = nP_216_216 ^ nC_216;
  assign out_S[217] = nP_217_217 ^ nC_217;
  assign out_S[218] = nP_218_218 ^ nC_218;
  assign out_S[219] = nP_219_219 ^ nC_219;
  assign out_S[220] = nP_220_220 ^ nC_220;
  assign out_S[221] = nP_221_221 ^ nC_221;
  assign out_S[222] = nP_222_222 ^ nC_222;
  assign out_S[223] = nP_223_223 ^ nC_223;
  assign out_S[224] = nP_224_224 ^ nC_224;
  assign out_S[225] = nP_225_225 ^ nC_225;
  assign out_S[226] = nP_226_226 ^ nC_226;
  assign out_S[227] = nP_227_227 ^ nC_227;
  assign out_S[228] = nP_228_228 ^ nC_228;
  assign out_S[229] = nP_229_229 ^ nC_229;
  assign out_S[230] = nP_230_230 ^ nC_230;
  assign out_S[231] = nP_231_231 ^ nC_231;
  assign out_S[232] = nP_232_232 ^ nC_232;
  assign out_S[233] = nP_233_233 ^ nC_233;
  assign out_S[234] = nP_234_234 ^ nC_234;
  assign out_S[235] = nP_235_235 ^ nC_235;
  assign out_S[236] = nP_236_236 ^ nC_236;
  assign out_S[237] = nP_237_237 ^ nC_237;
  assign out_S[238] = nP_238_238 ^ nC_238;
  assign out_S[239] = nP_239_239 ^ nC_239;
  assign out_S[240] = nP_240_240 ^ nC_240;
  assign out_S[241] = nP_241_241 ^ nC_241;
  assign out_S[242] = nP_242_242 ^ nC_242;
  assign out_S[243] = nP_243_243 ^ nC_243;
  assign out_S[244] = nP_244_244 ^ nC_244;
  assign out_S[245] = nP_245_245 ^ nC_245;
  assign out_S[246] = nP_246_246 ^ nC_246;
  assign out_S[247] = nP_247_247 ^ nC_247;
  assign out_S[248] = nP_248_248 ^ nC_248;
  assign out_S[249] = nP_249_249 ^ nC_249;
  assign out_S[250] = nP_250_250 ^ nC_250;
  assign out_S[251] = nP_251_251 ^ nC_251;
  assign out_S[252] = nP_252_252 ^ nC_252;
  assign out_S[253] = nP_253_253 ^ nC_253;
  assign out_S[254] = nP_254_254 ^ nC_254;
  assign out_S[255] = nP_255_255 ^ nC_255;
  assign out_CO = nG_255_0 | (nP_255_0 & in_CI);
endmodule

